`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZPVr6gPhgA50m5jEg/cloU5pPzs5ur+MQW36xOcR8MdF8wWaUr8zIKTkcmQ2+yydX1fZ4Dyi3sIY
TpR8Ac269Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
m4q9MtEWGVJ85SvGPq9Dz0jIl7zWLDc7qOxdMPlcTg9T1T9M5FPPiGgkxREX6nE7+9JKkFDwnsA9
8+fSm6Oi0bE3MkKI9FO2ZXM7K+4Rk8vDA92zhdLKaJ34nA7vjScrX2b/LBmzP8q6nQDO40WeaUg8
L807mVHk8Be+E1biF6U=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aatvZnYN0uh5k7QSlNnnB6bvhD3FbME0tc3JI5aMmMGgeBi70uOFdm+jeJ/aiZunLfXWyCxoMCdc
dBKB//l+xg2I91pEyCdzuoUrT048IsBLQwoZokH799mJgNx9daihUGv5ybbWk1i/wA12WcjDOJJC
Er52KQagyjyU7tEBN74=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dJns6s7QA8cdhO4jfiphF7PmkVvVC6Dhh0L6aFNskwPuc6Jos8rWXR3Jsgb9Qh/ak0KSbr9NkeLv
RgWhqRWe6LELfKQmcczmKfG1JTRag1Ex4E/VjixkGn64jC/UtyXNaVM5yfO4VMr/fepoyu097gcT
77pUFtteJrLFft6+LFiCSz1u1409YDqqA4/3ehiUO5JOTCVkxneqaqe+aoE9AvaxJhXMmJbXxuX2
8tKWpWklIhCC6AmEZ6vWD2uWzR5I+9OwtvmDMR4Kdzhy9mgzB/ud3Zwi7GCYMIYw3y7JpPsofCgb
v7QgaSwvHIaUuArSLJSXzaiJo+vv2cUDfF7Kbw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D2SIfMgicSOsDpsKHm+y5JCS0B9zepyfPIW5qstyEt9dSu53QxJ8dnCG/hq1rHPPNh7Ynj1WE5Vr
omRCeZE+4pAJd56hxgT6gDGsB9CWHv564ekGt+/ni622rk32WJgUuR1+z1V93RmKfyOTETzifJzW
c87TjOtsORPS4hAn8ZDvknAumyZPKMcIx2qqbUG6HkU0plfnmrKVtvmQFuscX/So3RuqQmaVrgEV
NxM86dJR4oU66dzjwOUynRyBsQ6WtLWtBkJ2Q58nTXYozeEQ2np76d0RpZpbLNyp0May2HmzXMGV
nCucai8VYz/d2AjP0bysze55WqGsL+qEO8jKzQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tMh7AxjNYMBJGMu4nT7+MUezQs9H8HlH2v9U7UVzGDM33uFa169W7t3PYXdwUnixdASrg4Ii+jDe
wcKq5RtvD55ebjKBFk+AJkdG5+4o0RsJmF8MRdgGUjYsu+yc0E70kG7GISyz5If8VZRuf5sfEebp
MAVhUoIklYMjXV0641B+WCQ851H+VAB7G65Z3dPbNwkIDySVa6ZdOY8Mh7SSRTyPs2u1iaLTACcr
cNLUc3i16RbKgf7QG7DMwDeInwsRMlfNO7eZeGEpaTeNPJNGd4TDVZJBkI1mLP8U6MFEOk+3GROr
H6jgeyhRsDgX3tTSgmba6DM90HFy2Y2meS+LLw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
3vFdmsGT7bywQxjNOo3Buo5RlQwrKqE+Ro65KpWn8LdEYl/GTrto4gQ1v66LuqP6EKUxiV/E6VBJ
k58NJlb3Dcf7JaUQhMOHagPhZO5lXenYpZxfscxZrqp4IweOdOWBv6vdozi/SXHot6eerezcK4eF
7N+40iwkuJyljv+FZsL8GhWSAgBEFyyekA2nZZP+ctUT8EkQ5gXYyzDKVjLNh1psIoFIQ0n1YoEo
oyERMU/yRCRHSLScNO9vZqn+ZAVoXeVZFEMV02Z/f3m+P9GiCvlpNxizICxZUOd7ZiRhhtQnn7jH
CvwkgBz+FyJoJWlovKdKgqKRP1eCdBn9dRJmzYaINODZY8kHD3+bHbX3EzUfkRyAHbDwW+4xHKGK
NJ2SKOepfMfhcq0fzeq7RIGg8M8REPgt88+PPhpFtrHEYcD/hYYpH/pjMZg09RZaGAnBcP1gKr+U
S9yp5qU7r5wPofz5D1FcEvTrzUtrVMBa9vwTX0+8SLgrFEiGU2q4eJpkuoS3m2ZNR083tflrvRD0
nCBK1c+ln7NL6jyVwh22Rf6KkSFgySBZtyIlyDtFr29RDo6mFPTrORxAh9TZ8ndto9Ylay5knYn3
3Pe1fBkXwFsizqKyg+KlK+qwHD4fpE/UENQZtaRbb/vn6vTX9qQG/SmORIO42TA+de/2cxCYft0k
g94biGumCue6VaYEPD/dWfC6B61SeG/CJxoJRan1EWR1GvqAv22zF89cO6+SP2p1sSDiflSywrWG
n3lC46k6Wsw4pzc9qCwQEEaBEHE9VjhcPTh1IBwFr5NaE946rzOax/G94yCY2g/NrkM9agdh4j7Z
P3vcDDynkY4fVRKxaJWF3/5dG8sw4vSRbdVQJH3zVjaGlswjDieXlzkHPruup2x/JPe6zsF6eS1w
RG8CURP392eyvU2Yh0Qy4yDiUibWCmUzsU04f5JKCyzazPlnbpS/Te2CeS+vj6SiX5+2K5mry5aM
tGrgDuaoSl8Q5dHG+ZKtIS7jaYVnQzVRuBgo63BNdDlCNXu6jXWRdNbKuw/4gSxyewLYO/W9nM/Z
LQd1bJN0xqQ9hpAS1+jN83ZD3zYjM/PgGz5VZzKosJbKhoItuW1roBrDQi0K3OLuObisJcjBs0O7
Nh/MbIkJofxyP6rZcNDQvdYs5jlm/uKf/dFQQgZE34n6wAZ0obxyjTAPcG7dkH5RDP4o66+HDrHF
TmJ0nN+sr/qyBZUTIym/i9+YcOuH309G7lQEUDSdG7hDdNPPJmWBNDTFx8y4SZC7t57BceSOdkC7
Ss7zCf6ONWs5GM/AWFpwlqr65zrmHJoYuB8Ri4jJnNTATaa40SPyD6BvDUkX0MQdAbuIx2evaOUR
2+LmJUsLFEwdbkYuj4425ZtXf/YUxw5KHk4q36FEXntFoXDl+2ViZSgjRPdkmLpE98j6VdVzpCz3
VLP708A+CeQRFAGgQpqMIAjcpcGEIYCd7JDfCz5dnaEEQjln+84M25rtvByRtpY0xvVL1xujwI7Z
SJYRiZKaNKF0QxcPNKBylxGD2fTp9VHzy9NYCNyIvuWxKl2DRpTqDLI8jJfMkWu/b6rAI9NoDRVS
lAN0+FGRKo57oAdt+s9XVALkZ1QznbokIm1eKZh1Z1C7cxEBWjAnKEDuMu8WfKxX9G1ZTn79zt8q
8/UOEbvZ5kqCYGdozPVqZZXXC6jNUoPDH4KeatvJkuWRLk9vE8KW6jCabo05741cWJzx7XJXL+DT
/Xq7RcKKFUOS2yVnNP/oULxeROHgPYH9ev6Jn4FrHHpwyfaY1PvOhXcGVS+VI4xASsZiZzYY182P
VRTfFT0cDORnkIBdXVXUbrITsDIcltOp0sLEoF5eAmLHhdlpwBtwSfjtqdKUESTVBPkbYIJH9wMn
vV/CxhDIdAoXbXWyhqOxYwbXIzz1fIgX+LwpKBcFTRI5V57EPm33Xh9udT5eP8MNuQEqgzunLqHE
gWAZumXh28diDFcsamFMsqi7FSh0bxdTi9P7h7IN+kQG+NtRBStHcbx4H2SeHjsUK5sAH8SOYtta
pox9MMuHG8tb7sxabmaXpVNhNTc5224JbSJLzHyjc31/GVLX2AZ5VLRByoNQYpLud+OcqXAWYHLo
p7FmOG6krZ/9YLOGHfsgn+nei1ViDO8o4b3bhyjcucC5ZM0X2HBjSMwdmVNs7Ewi+a3kElLOHcBx
s3aQkZ+GaXuJLsmBjUUGSPehnXl42pS2MeHJxuE7J8TaEJDIDmuvP/4Cvkju13OaH56IuOJYrzD2
NcBmm2L5G3nY1ARXCyp05DjCfbrwNqIDI9iZ4eQ5mNIQD6GBy80AtoCpQlgI8j0OrLM61anygZ1g
k/F3z/HWJuU6iTg4XbgsTz6sCqkVQegnysscsXmGw69qJAB9LmLusL8ylsT7gcOFEH+e7jq41OCh
du4qzmGfjVQf3Ky0YIhfTSx7UqR8tMVEBzk5TJwryysgwft+7S9VVZzklwy8u5UxxfPTZhS+6tCH
F/Il3ydBdCWqm1XuJ34d8zS7F4gCMQVGTOh3Fd2FCuja9KQa7dbkGo7/iDLEhZ7CS0OdjgkSwqMQ
YOQZhwBv8I8pYFfC4Rfm4uSwCHQ6/88ZNFUdA64AxLgErMLcvE0vEMP9UhUCU4vugfFCmiDBCpio
2/ukfitOlivpavOFT3yWu0yhcObg4kS7lnS5jkzDmHMMDf2m57AcEkfLwTQbPVbUxG6zj+9ddBQm
yzUZwf5/C6cj7ovKG/5z3qhPg/1HHKsg26jK9UIlFH4w7odXi89CKR5/MNHiq8dpePEcLYZeF5cw
qa6vkoxXjp7lvmpwO/nXK1xVDgLR7kafqigogzorqjuAdeTsU/ekdWQVP/n4lwbMP8gvSZvoCpyE
zF/E/0gzBr3QJNlxCxT7woH55ai9JV2X3ML3vUqHP5rp2pRT1wHmB5HjGc3T6zTObab+UCx1RDN2
mzmlcf01FSS2TFoUCYPZhiuOMc6M37BcdFUZ2teJoiAdH2y0b4dIAYlraJ5uYp5PMCD/Tms/RfId
S1vQAzpc2qGlfIiOCSp1r1P6A73Iu6HkY8sphB6fbgrUubdG09UNcWtevtA5mfTkpo1pOCYrNgls
atCU6/CdLEno+Z4YPxLdT5FV4KQWc2zQiWHWqjp9xTSycfUA8s3uBpCr96tcIlpSOunLDHo48w49
c340iLuqUE1JlIA+44yRsHizeSKHByJNPQvPPD/qBzf9xAq/agpqALGCc6jx6E2qEfJQltcZO+IA
idlyMlKVkhQXTFola7nkx61EEqT8TRSlATn2ooudoO8VEfkt7t3IfgV6wuwaw7bAbcJlHUnj6sH5
X/jtLMA0S1/rOWeVm3R7kv9gamXQxV1doLfvr9+rcRoTGQoICjonDk3btnVACIsmxl1NRTQTw9Sr
adC3LiJoHMifQNEkV0fSXvPuGPATODihiEJ/XwwTZt8jT7xZ4VKY6ZPjRHmjojFT6l+YL6ep7fz1
MVDXsTEcD/JELzDo6cnYHVQItfXzgwsfZeTYDp9O2yNtv+mJQRJeHll6oEKrhi62zzwNE/EZujhL
18Tmw5UI/wHhebVLaWgLMuZM69d4ayLUJ+hc6cy1BSbHEG6UnxEwoZEbBmpC/ryxsPjhxkacTvbr
Lm4jDnJvJAfmiCqsbE0WtX1CCwKolnuIgw4MtX13xOaGcYRL/ClU+Hf6bx9LA4nIageOwjREx9OD
tNO5ryrRcYSrmlIXGTeVIBrZxjT2j+nn3BI0mPfRXNSEatsLbOEjKe7s+Gh5N23vVZVjfrPF+D2g
fSVHScTMsOlZLHFoBqzk4ogWhvojX/fqwWep/DKh7v3Na4u6SWF+wBao3AosWpG8ETWCuUrRc/eC
fHafmIwPSEZwn/J9S8FjiiFFJxrdxp5r0eFzWxGY32AL0q5LOkuNYWKru5f3L2i2ir1z9iZLeTXU
UQ5/MdbjJh9gv4W6kVuOXg92T6MvShiO8m7+eCECVXax1CmwlpQa7Drig2XRoxSqf7tLxi+jXhOZ
ai1KefECmr6BcqQQfRMX//D+IicjQdsRLtes79ES+R9NZTcfMOsQrzHK/xZEbJgmIPSHXzuCGyKw
U31TcFh9QUdQH9KXqOk4Jg1REKQvv0iYHBY36x2hchmylom9vvP2G/CDUcgh8SRx8m7NQ2AXFxrD
HxxXr+z5sxiPsz4MJR9GA0OIv1UW9CVGrQPHTjzyt8eH82YEXHL1/lLzYGVRymrr/c8uJ+Ed54fi
lLwbkutDVUspxCm90jmU7gBwxZE+7yGVlJSJtqzS7dRjG5UK/brUfftYHjx+hJpmR+r4Ja4GmZUZ
yYwDpXeof7a4B+lMImnWpkWUI2a7XBov8Cvb5EbBkPBqRa8q4RsB+5+c05x3dxBi5r+fVOa9p82x
p2dPcyDI/A1dwD/jZKElyMxst0oIYg1G/ZHvgjqUgYCSRUl6JT7YodML+V0WH+n6kvX+T9wLveS5
Mq2K2rJ+09U3I4kRUYJkrGxgIuHbQHfhPYgXv7qJfhLMUXdvbbr11Jwee9BTMQ14OoWXrfhU467p
osQOL68FBp2aGlOi10BhJUopZeu9aFZQYF2hEgJkowsx4bgFhin+p/eLimX5dYMRTV0L50RSmfJ4
Phbu077zJfuf925x0vIZGYvf93HO+C9qSlcujhPH8sltTqOIAjQoreMm/Oci46XPUN4lJGGzKnlE
BtwgRcYiIcQ6Ph/HZxoOwvm2OVfWkxoIf8YBQGgHFi59F7q8oMQ6sGlMvQURxcxS3z+MnvhSULU5
oWV6n6ACsnVpMZaMTYD5lLzerniRH77RWWX5QGbt1UgdzgDXivkfdI9Uu6gxyCVUolTqpeyaBvJU
prHEOSLnciclBon5FWSONB56SYLH7HLmZVbHlsUqlLKnsja4E3mgpMhhqQ++yejw5MXECrSmLb4g
6UMKB2HtYHrP2fvkWdr33uVHyER5zFWKmcjpbPHbqlSVF6FMFQ+TZqvpnZhwYZTUXC0P6tCL/jv7
PeBjIAUwBY7+Q40XVy5QD3yuKhSsDsnAOCMH06nomitWpUj41d5M0pH2Z/dWcJ+xfcilY3Q0Tl3p
BDar3jPYRuuZ5hAGk4tVyU2OslGPC5tb4lmAyrGo5AZyi+sLF/tRPhnzA2DOqjZSqHVitmymH/Ig
VN/Pbc7nOCTDZ7fIM1iagiyoFp0y9YHeaer5oXfx8tJecpQte7gM6nvffPbOCcKM+N2rz0BdIkYJ
mt8M8b1gUNT5eVg8uZj83iN67BEput/3IS6+5tXGqESj74PsrHwVw+iP/PqC9QIAuQMRBBp4I1TV
iFUThSgobIe6GEVt+C9Ards+WHrQJog3omp0iJDcCE5FqkjVDnP3hPi1WMNslSCLtaYuyRbL/oyu
JAzhPTlJ0k0drtkpO+rjd7NkMvJ3Tlp1oj40n6sGYIFWN8NTw3K5KjnxvVdz8aXFSyZXchwWKm9K
t1CZZ5D6273PKuxMdUAEdkMeV4LoNiz8Wcifha/bjgXnFjAygOF5966j52+Xy+pzfYpMS1EziKjn
+IXZpYGLjXXHIVEBT8wnokgF95sg75Bs7zbFBlu6qpJIGureEOGAgiX3yefKXI1DmanqqMRVPJMu
52HriiJntlibUuEHdf6qpyxiheHeNHfnBUWEVmIJewuNeAqosGUGpBuX/fU4jYHcZliRLXM3lvf3
krwpNe7NyzIvSQe8nBZroppCvw1FXscP3htE3ufIfDpQceag/CllA0/d54WWo/hM5hsdjD38lvxn
mpR35jkmAsOP8GwbNIzIXjZ9OYe3JxmJ/5yuk6xiSgazIH7RjLDDQTuRPvGSXTP2yN67flOz6zwc
+GGnHr/AsC/TXPvnY8YeL+Qi43OnGWrwt7kODDG5hc1u6ZllB93/3nRWQKgq7RvXxTjJhmSoeNbr
C/y4fgEnBaJDMvAEzoHvtcWnVezENLkzyr4hjdppTqjCCuep4WFYSTTbDCT6fj64Bt36KESP0MXu
IidftfvQQLf2RcFEoeD0GaEng19oJ3fyYvpJJntF0G48oAvPjyPAEDWr/PUwKGuXfsRdw9Q3OFAQ
CURrnGCzA7SzukEwm2xZzUmfGRrRca+0aIV1oC4Z7THXfGdjruWZTadmPi45ZDZrZqtwUyd/yiUj
INeIIWrIv6rAsCQwIZmpGWtt9/IMJKUyilclpG1vdcvXck1PKPMExcEffGY0Miu6wM7jnusLs5kK
veQlv3+pgNBVmtDFf6ZEXQeWD1cUkizXplsjR03b2l8iXtK+F1tcDKhMnDZt9BAe957Ukob7nqMF
uQ2K/PkowZhIp65nAh07Rc6LB2D/QDfSTwIpuBiZLo51AVOgwNJIN5zvZcMYyqxq0a39cTWy+mvj
jlLVSTnWe2nwNDUs0miaacp7X4yNUdPaq95GBPQDRGAy3nx5XLajgZLjBX2m3o40D5wREZxLB5Dt
mtx9VSnx+16a45d9Cch/mKhG8CUPrES3evhkhHtq3vCWmuBPdbb/0RVkC/Z2r270o5VlmnZQnLov
QKq01EGP1vqdKMVZY/e7vY1YQwlkBiGwXQEMiOgMGkXPCh4mqCUPp57NqDheP+WKvQfrQPb16m4b
ij43OtNiX1lSPcLE4M6YLSQt4stC9C9+Pw3rSyaei/kiKHZMdwz2lOCmfL33qmnUX/yj4SiCTmBA
Ka87ERFlt2jYOgP0dwMlMgZ7E08iR/oZYdId2wrMDY4Og+9LGUiBikLY0i8m8a+zqQAObiBhgNaA
wMJ+AWaO/iWErHJKf1Jb/PX65gAO+gP2Ry0DwerFCSANy0R5p8Mh2tF7Q4avpTK01FrrlZFKwzJ+
q+X1S2qsn5XGCVXEbjkxUjV0/K1RCzBxdNd8iUKJ3B+0aUeZbL/aC6Br4p41UsJKAM9M3XDGmYZQ
75fA4UPhRvpEAjbunkuKzz+zxXAtZw0TbUNgO99Rg10FYlp2dz0Enj2IiPiCABce28kjPR5+9PGF
KL1+KMZXkkc8neW5w/rGeOVhcMlP6+oEZvLGgrjf7OwQz3zZXtzMa/1M7BD76qJwLzpF/trD+xSL
rzwZcRPuAimKm/flPQCbS/oeWXD14B6eq8T58McceSUSDOZOo9GGnuQWskM2XW9zu741xHeX/85P
r7LzCCjTOQaTZzQ9c5yqRYKlnCH2OGdzbPMqBarMaNaA1pCswij7RKb4NDn2+B29PQq7ZASa9DyL
PXdpy4Wb+2QnmG9Z//V6uGhYyVX6eF2EzwuBB6g7bVPret+0/82vG6BMiHzWAtIpc7Iq45mXbYOu
9Kaf1hMRTr+WilQGpgw6+yCKZHU/wwn1elyqMPEykN1AIyu51P27xC2MWcPGDeeBOV+W9BQ2MSvO
cxz4RmPgu5Kba2IvGoS5NFPiabKZVbHxXkIs7Dxcn2nVeWRDrhr6/V+7qIAn1qBOIN/bADhNEYY8
9jPZQTEHBRHGX80IV+RamN9evzBDIwd4EBYXrh0QY798Yy8Zq1BmeO7u6bW08e2/r3icI3xsH9pw
JC7mg7WtYOb6mSWk0XSZqP9Z5PFKwtcQOUEUULjgUwwKa3jaQoLRMpsFvGJYJJArq1wj6MTTeVkt
F+qYlvwooxeM610AoNyJIqfmBlYCWyHLkpaTI533nqi/lqRpXQvwJz6ZGs1LbCODjWqbYu5ql++i
obhIkFAA5IAXokpEJr9bEZ90jML+mHI8XJ7R/SmN49V45jZ5I7fDGvn/6jgLeSOODjd7flq3C0Cp
Qsrxih1qpfMsAVEGY1rZo3vZw3FYQU2kflRipcIswbAFZKO0iLTgFSQUe+FmmBdzbMZql555oOnT
89KAhMkIMdEXtowDEj1IS990NZokPYjVbCQszoAKtANf87f0ao7cn62cazWFEF3bB0XCP2kyzVGM
eNzaB41lohk1s+F8g0KMZ3PwczjQ6IdcC97ycl1fP8PheSEYh3zmth+x4U/Mv3QEnbn08or7g0TG
P7sKpf2SYROj5mH4FLilHlkFt/2aizkodC2Lla2bpIYleKULMAMZrQMGeREZHs3Q8mcLoIOPXeEq
mRy+bT4CRLPDAyc5c/YNSWfkscs+7tPhsL1g7ZxTEM19VYNBEJTld7LA+1Jo16pHmm0lSQ1rHw14
luiELmqvTnPJzDMMSGxdLscHa+RGJz6UPp9TaMVDI49qRuhsPo9Opj6EgeW6zINRF51TNyTllLge
gAb7oc0nAD8cNU/oOd2SpY4x7BZoOq33o47zvySjVLf7eMgy3Vi91u/0hYm/Gf9fHodHWQsrVhKg
UTurlN3toYrfAgucs0a3Q99xsy7FRe0qimMkEoQHbhpCpQIEV8JocGI9NCtoAn3wvOYm1a8ixkEe
jg6tzGqvJ0AOADqQS8tAy43DCU01dG76HB4GE+g0bH1TGoAo8pVM9VFty77te2GlkyHyY+zNmYss
ZOEd0asm4oC4NoKKiR/i5o+cvzzEQMFA07bI0Q92helEr7sy0XeZzdjOUFEZYPHOSgkqZ8tVJzIr
fxDKGj2spmER4R1/AbSKezLMmxpftC1wPQTiDB+97CT2U0yvXTB7fKLe8nehu3eB/vBPtVtAAGz2
LffDJXb/vuZw+IvTc+FC/UFyBcW8j59KWmBjTn76uPviIXXlw/q+v/e7JYll+ULy/PT8/8fhgjG7
d+uWc6jYE4G5WDEVIqxzt3tWgiQc5zYmLeByCXphb0pLuUcV/vKDuF2Ro0cpx77xQTYCJHDGSG02
T+7g/C8bu+03+CzrOGeOwssrdJBcu0a3ZmyBN6yeaB5y7ZwD+UBMFoupBRzYKP8w3eMVmQLmR7dx
1ggGRTwsrOGK0WtVgnzA2Rc222R5eOFW7mznsqzkOqPMLJ3XHLEINLmCrtZeftLBruSnPaJv0/R2
TlTSeQCEUtK5LJYnitM3XvSSHMPJv4GRuEbZ2tF8hC8BIixvnL8F20/wMlRXPYlcjSjpBFWLXEk5
pddSSkmhLdfnO1S0/g2YTV8eLKNeICFdPyoSIlRcpx2fMx5rTRbIAku3YpXjqWGGQiueoDc535gW
/MYhGiomXCBmnvy8ry8pBQYYE77RdLE0Mbbp23lu8ttD6/c9WhXlonuFbnPX03OnA+SYxPtQRSuF
+SSLFKOosnHnGK+XL30vPpm+RfK/a1eRMLcRt+joEaerzlvVCRv/6UIYLO55D1jH3/hpX0eyBE5N
3drJ6BhGlHTG0TrsoBiCabn8/KCPJW8U7XsQU+D+qxcsa/Rp7ovAjG/7+Iyv0I86eGXvxyJtgwiG
Jti4pDzpx64BxEGFgA5+QdRsW7Wr4pUFyWdctwNxnVVp2FBbU1F9cz0NW2A243E1F9bU05uvSBsq
7bJs3d+O8XHcG0fbTgjcar22UgYL7i8EaUzGFnCXup2QbS7mdSrr51q+G6nBz8MrYGB2OGGvJwXM
VkscIOzr3RTsDukDzpbHcoV42s+iAmnQf0/sP2iMTQe8mcahIV0Y39GDqUxni4eiiCn0kid2fRhG
t0GQfp7Pqh8CERu1Bb7wHtYlvlae+knNLxhSCOm5KBbFXtfO/1SSkxFWyZ7NDg3UGYWNN3/pEwm1
eyygmXdr/NcexJqqs7PfhgSd8SU15rgnzsdMAF0PXsK6oVgTm8V6lIkvPjhD9llgvTYHRO/bqCpc
TiGNSlAq3rAb+LKIPDEwJc+GImqvCwKwQHHzJFtL9GJCmUiYPbLq3hQjhyb+vGOamfkdxml6p8Yd
owZuj0rw48BQ5Y51G8xkEh40oqL4YtzdQavAKf7R/jEJduPDhgtAx1kftZTOP5w2zFAaDzL7bBrf
gsbiJXcoB8n7KiTwU6gzeOrQsTiCPFuCE/v2sLXx9Nny+l+K0+Gyvnvzyh66pj69yuWuiG2uitUD
5qLsxK21FVO1oDSgB2vHG0KZdMfA21Is4dhSebvtgkR2kKLN3koOMeqUatGL03G6zUCtkn2IBFzz
JsvHPkRIz66cR/Jf4Qr3byPXlpWQB8FO6hD5krAPtJrlaROMWzk5o8s9rDwJXdrY3xLdlj8+9SHt
En+vZBAbvomzrlcE7y8GF/w4sdJg8Z+qN0hmWnjlZjvz+UCHMdtUj35919f2DAVwfGN+OxemGgfR
vipg9VCakdcHiu0QXMT/LVSbBjs3CSb9zSbZZohxiA9HJQponuzKVVhLxnfTpZUehpsLKCTXL0vI
wMYw9rSLYZSF/bWLgvZOy3g2e6fPtOl+jtAIzzwe43MwUjV5y/KVcqgRB8+ccUxloLXXWEdd4UX4
4PxDkZKpDHRbbDCop1q9UYNMWUtTwDHrTIl1ECD2RPFDAFfa/QC1+Th6nO/rjfXZLEboaz5xXIpP
3UIVqXGSnRgHLQ0MUczrXIGcPEQMK//n3UUQOndCozKY1QEYgeFsxa9DPIsbpK4PDteA1sPfyi5s
D+UlF03W+/wG9tMbWcMDOUac7/yW5+eL+X0JRhQxv+pD9U727rWrKTJfAV4PJy6Rg20Zi5kiLKqC
ru+9rXtPl9723qzAnX1a8KrHA5Xw5gAEh2Lj9AVRUoUI1UJme76UdhDhh0Awmy9d3dEfAtOJLnin
IW5t1oEU8qGVN/6V8/epNZLANiK0YGTtTsDFRP3zrXloOor6Tpr9eIK6hyy49RLnwWF/LriCbAr1
G8ZxRSWN0J5TVg+VKaa+xdC4Mf50Q6oHSUFMXhfVCu9lSGh5/qqyHYT3SaPN7D7NakpwVpRhWdfS
5DaIMvZaOfvDq5k5+gz1muWkW2xh5RJjegAnH2zHfyg8DhiKRPhdtYgFhUdWkJ3NOmLY4u3AEDxa
uzVkKPbUdqXRZNAQyzmFATWifTH7eM5mmL7TVRuYlonp42KmOWrtAkH3NzgcL6qCBgDIwy+PMuRE
FUzzYQVTDMIHYtwzAc64k8wc8OTolatYehLXFPFhJadCUQmeM7mLAl1xqABfV2De40SZbF+zIClV
cADmElJYoraLKpSgDWp3Vdge3uxt8UznoZv8N4yYHg0kiP613Dn77R9FJ+z4P263OvWtUSWVsVEH
xJSqz8lFRLFPRp+kf5ZW07Eqn2fSXqRfcelsChbE2OZfGsv1Bo4R0bpGWvFpbrS+NgkY6WmdVeAx
EfSHR0CHhlenC5/FBic9pMQ38dWw/GD3UC2mc+P9p9/DqYrP6rZvPxtJlWNDsXYptgFEauBnFcvP
K4WCKkzRH1OVbDMuvN22Hzo+V6Teki17DHNpluJqXal3DEfXkswsY5Y3eMKEsXV/oxiMDY9Coq5V
ws/7IepdBzvhEcI6gG+x8xkkp6OvGiu7P0txMVqJowUOFT2MCyl8JIlX3fBFBkgaUxRk49OhnW15
97KAnUjb38mUte1d+SoUEzOGZvS1e0sUmWkpadaIBq5/QE1Nbx9B5dBGnZl5p+7eQXe3myeYsAmy
1qURoxTwZAL9PasLlOUVbqBxZoROca//QZHyEM71EJchVq9Ge/VsopPtfsFg62qKSkSirNeO/lZQ
smep4mUVnqdkKhPsuU5WB4kGhPRZWeaGNdLBWfYQdjZBSVumSb4ZV9S395fPsVbxSzAiqTzqHCZD
khIr+WKMBaO/nC16zn+9T4guF4/hK+dima8eu4gA4UDAZgESFrwLt8q0y4wsNRUjJ9s48UYrwoJS
IUInIY7o7VR2rPsSKtOKK6mTqpZ2xVjVaQ9pAVCDUa2D4gUXNzReegxJUcvkLun6/yjcpAEpn8zh
fwDv8KlBbf4rpabtmcN8I5MK3OnAskRE4mL8JUj343JRfKhMnCNgu3RlAQzyZ3g/tDgFXY8bYlUI
fgSNyL60wYeAv4J8yCffFNIzSNAX1qFPMv+iEiwLnhQu/6v9gqOR5lcW31SSFlhd7upY/OpIxXi7
o6hP8uWLOLhrGYY+wuS7Fb94NHCakrkoQJk+j9+9bEk+i5Yd9uWA5ADUIFp7J9e4igWh4akSZE5b
L6h1I/oDBqah/XGrv9+25qnnoi5E/ajMhrFaMB/toxx8IIYSMTM+FdipmJAADCNT2YDgdffmIJk9
6ECtJhBMNFnuOgPQ7R871RAcrXDFmNB1NOmNq1bdxFv10ueXmTiGcift44gE23Y3SfZ2vqbve+dr
3xt+iW6rKJFxT2V1Uls2VIkUptN4JzxsFwOpaLCwnDcv1RUM17hSjansltrC+ts3x4w5T8KRFXIN
YLVuj2Jdp05N7WZxdY745dw4fCetuKmJv/mjE1omQesqBDs6o/vhmi3EyKjTfnY9cNvJ9pD0V1ME
yRI6O0MNOeDtDWmp/BqODO9Qsf0XusCgS2+YLTZZZd6ZNhw7WYzwjBoRU6HuIPH3DJHX6hYJvFF3
sHmBpRnkRt4lAKZ1ukpNxbuMrTBE2aM3qc0hZE5vsLZ4C0PkejbGnpGRvStluqOkJ8ZMToX8Xbkr
iNJuZjDXlgKAkgWrt/AhguvSW0vPc9ZDLSrlWxvh26iGTcteUu8OR5uA3g8+YTaq8mEawrP+wgS8
f6n/xDTDZ5KB8wKI5b71PWjDnjrKB/ekavROfbL0ee+BAuoFLf+ts1LdwR2lAf44Q0MXWNB1vTnP
Bk3lzIxUY0bnd31g6Ys4uN38qro0bAw4+UI6cJE44xXo6pEMmbl6CtFBf3t8jDBjf8973JZn2quq
7HlsTYgx/xreSi9ZWqL/5PXMN7VIi03tNq/TPMX70rGWXrItIOWMUPImlViKusZpdONWzWCd7EQI
RSKjfgvpiRLekHd9XhlKj/e6mEd1k1PzAcpvuoKd2ududL7WBKVMYKdmxjfSEs5sg1wRPTY0xBDb
7aknHjmEYsJTTcsrnw6lLrWZcVy29t9Flco6E36LD1vrZ6vdM/vnbaUoE2GMgr7QjX85wnK20eeF
21XtDwayktByh4ncN2K5e+E/ziNefsUx8/QZhZtBcLVzu+5Tm+gnRrODrgHNcxoNMmkXBBFG/SaE
niS+DNTrrvRbADso5t1nrcPo2enVOe3646hiw1pE7hdZb6uraZKICL/AVHWqrMEZOD/KAlRAhgIt
8gyq0g9r3NsMzo8Q1hOFMg+oUyzyOEU8Q7LWTOXLX0tav1mEJcutArv4P2OWGShqEYYYif5wPsHy
eFkyZAqt7YhsPDDP21yIacMLfy0wSxupYq8yRjhiHZk2E0R86eA3X5I2An/1E8V68ySFbFpL/BnC
+vdnDO12BJ0fRJUmp2cA1mRtHTmXVDxh7sk+yfvZySi5uXAA0k3+2kzs7Q6YFyi9hCr/OvjDbXGa
mV2Y5gqNsMHHKPyAKl2UfTBAV8lMYWYhozcfhRRMFfkA7zVyeuJ1+x26N8cjNbjlL1/WHjw56nUH
MJ63cJEra4UhPbrEeZxP8+tM4vq/9mzOaBWI+GgW8C6zKw/Wd9YhT5FPHkLAGrAkdxT6RXPpyPqN
iXcXK1Ls7sX+1emmX9SYruUcbAf3Qz3/O8bcqdTp/fyMT4r8o3We8t8P69+JlN5J0ZDuJdloAcRI
uVAovi8/rU54TG+BWnNVO5Wtq60pArsSRzlC47tJpAW6IAUAU7yhuX1oP9RqMr2EIWhl53RLb5/H
cHdjUCLuevS+u8k9RTDe6uDFAo1msYDidxwcsyKv+a35DjnlCuxOBt2QTKcSaooHUw284ib3FfML
Im00nNRh467NLx+Z5z1iOQmsEzxAwk+zU5kLinXCZdXhXPd9lU9aXxaQTyqzIR25QLMAmZRnvGs1
ZMGqHqMR/kHJZ9WEQy2XVw3y0GcT4Az+5zkY1PKT7rA8G9fN2s1mMOHHJqPlkVDOB0lCaZmyRvPz
w6vgxKcjm/7NbrUtLLMEr/P7E6gObdKbQCiog26wZi1/CcbjBbfJUAReV9wumIJjtS7vQzqtfShI
v7rSrS0f1SIze98rOxJAoiGCFJGvwF4vtzTtRkHey00crNNX4jLDsXdZ6v7OX7uWvHCjkH3277T8
u4K53oNXg46IXT5uFinplOBV6GKQ1wfbfDU16VIR/Qoi4ECZL+S7PCOHzvMlCM97jrqqfDBsqLTB
ZsQqLE9KpWLhzBIXPYGR9xTrGHA/3ItS47YYGuexGfzeG1Hd+J1kSsKcrHZtdBjRg19wRugV3bSC
2VBXVyqtA96tzE3aKmasDkwlFB/5r7SRg4p0Q/lr8UK0+LSIuAzQy2CqE56LR3BA7YtsY3Y6cbU/
bRGe1YmE1R1MnLECXh5qlLlVVx7Vszcnpu4dT4oWh7Flx3ZaJZMPwnXpG+Om6TdtdJVEtRaPcXLv
7opbYYOVGe94Tv4o5NCty+0C3JuT0XUKuf5P/CLXTS/71OyxaZE2sTDO3MDx7p2kRVsvn62WxpOS
MIZ8dQHyVFgbLKTa6moaz3vnmb5pGwnXXUgc/QSo/4SKLG6Nj9EJRWNdW18buhDTHv51MJSnVhea
6Waj8xHRC7se3s9nWJ/1RARuBO+D8X1eL7tQo1hz35xgyrC1dyaSNv5F7XoImKf1TIpUM+sbAwHV
MQ4+hxjZoIvlulhzXzHcoLPD8+0pv1ZMf9euTM8aOBCLumicHtXBuXXHjFcWdd4WSOpJmCJEp00W
Gq24rj3mml+QxvvoNecI6sWU6Z/nARNo5O0vb8jDwM1p+BM2iaSgHh6ioxlBceG+JIDxGVFSLP96
6/kIx0rBIW9lEr/3jea2GeZ8f4xWfaFtHFip24ERt8hwezihAy/wd3+ZoE4oMvQddYEDDHBGv5iE
i+WSZ8J7vQKMZyv2RvBiQ2Dgwhdbvdyf90VjoThMjPvRgsODtE1hl1Pqc1yx7kItImJf7PyVjDlu
zMcHzU+HxPgqdL95SUBaseskuDOmx5DIJPAiO0HOwFuftQ2SyHoFYppGt9BD2cdy47KsDAhEq6aA
43Frx3e8NUcHelvyu7m2T7iFhoohWwLNWWiSuurEjjVrGZiEvNeDJWyB4nbpT+xlwrodGQxR08in
wN+3ESb/VfjJjx+myb3As64z/UOjNOZ8sMP4EgU778xkkNHJpaoNepE5fL5T65XiZ1G8duPzE2qA
xcyjWu42sp6C9rGY69Q+LJjOrgFKECiCOSYKH4ozc/6Ha/ijVKCmkREFHo+QLNtLMva1fclGn4HB
8R79iPSK1Stq2Tz6up6cOIgoDksfsJjC39ovF9ks38KBd4IsQF4DSh+jftDiC/+/MQbP0Vdx4KPs
Bl7HnvQbBpEHeaLmuPFA28XKgO47s+vhc/R/7cUeXk6B9u5CidaOYNVc7Ua2yuVghEAcekQAVkrF
1Wd+94KoCzGJFECIHDZn5Y035x+0EGKByIp9OmSSuoS6AVLTJnJOm5fo6woaQwY7uW20WhaP/aMJ
niSwGfsLGDFw3NkZ2YisKfg9uiMPTu9bHIuw3M97wireweR9/l+docMA459e6l9zPWN8yA+qf0u4
3yCriv8m+Dl/D/7UFM2hhJm+DgjtrrmVh7vO2wI4L9sUhYyWMvDQPBLX3XOF/BuRoxDCysCgb0DL
tmxJVSaB3ayzbAoClFNJOYf4DBvA91XRVVclBRa5aftfG4QU+ZPH+ALH9BXdsWYxJsHRUClaQ0uB
WTL/6rh/RjDt/fDzlbX1Q0EWPZQ5hubg7xVrr7tmNf3irA2XzRCNY7h3dMKhQH/drU/VqJ2jWtKw
EhsLBEtVQsvkaAS3eJOfBAXMMNwGeQNLweNymaRjs8t8z9eBN9nzLvnn++ceSzEFG0+h3W+Oqgwj
2TQHIJm7oAQ0dOpBUizW5AdpKK998WVj5F/FomWxYpLQEfgqYaVbYo0wjGVIM78JzHTX9By3Tuij
WXymKvEQBtt5GfIsqLSnZ3e/OIAgUqoN23JBEvlUr5tqIkm3EVwiHywzyoguHorbEHChd6Q9f1u4
WhKppFyOvWqy32M289T5bCX0+bisqEFHPrEDixtIdupIjhCezvMigbmFknlkZeZ4uq1t0OF3W0md
YtdHEwI8rF1l2weoxzoTdNQ0+g33GL2DC2RBShrgZzD9rKgPw7RR3tFpKwQ0gSkTawczup+Z6azv
y4Ukryo3jrTJd0Hq58Yw7fj+wKoWx3IjamSR525i6l6tSu5NEgh2ChgE1XgSj5flDFnd+RQ4+fiZ
VKCRzHr2oIC4ZkcJ1WZ46GkKN8CryDC3pUhxNJiNuo35007j0zLqjMlcihyCDdfEVLhZifgFoAHk
TiH0eZnBv+Q0Z8iF2A1lAmx3RHfZ+EktiZp+UAJ6u44ZdoDWHNgPJrrHReKRfYXXcluMF66gNZDF
lrlp6jNeDmsq6lhV5lkgzPvqlprNT5yUIDfW+EJ4Uf6seOgCiHcy0T5/v1x4YUK50pKjx9ytoSCY
UlWMKbxpq9CP6AA2bL/Uq9lnA6MYGYJxtI094m4QpAS4u73mtlvD0FqtVku/mhJexZirrqunNbji
AZiS3TdTB0mRQFQDxwiuJsvI97kuCT6o4rrmhvhvtJRdYVjLWCOHJH3vNLoYB7zu3TyVYkj0NHUz
cj6h00bxpl8MNwHXP81LMlDGLYT2NxgUQdncww8rbElVR0153A7eOiGzuKoEF9MUY4ihpVQjP2TX
4FMiHc7xgvYka5IkNlGT2BBMNN63YmekzEnRfmWMI8JjZ+fALTolHn9pdpLC5o2WJ2RLkdq3msRw
mQ+PeolIIIqWHTCRMEdYguftUFXt1ZWKItGTgAnX9zTp/TJ0ZdoysZAJPLSRUSFQGuuYIoea6/Mh
fxLzSLFJRndXq6vjt0Uu0FXACoOrFwzWyC82glRia3EPrL1W8c0OnvzhPQm6uNBhhrn7T+hcO0RQ
kUXxVZqKwZdJ7LPMSAs8dGrXFIkBHoZjdeUeau3uBLe1UUCsZRLZUwi/iFUZcnV+YrmdWbsQNevV
JoqBO2D721CByzo30XP52kaS4JFHT7fTmupFeF066+/rRN597QA04mBdSHGsDNWpzBi5+zqyz6Jm
08FPC+Mb9xiLXfSTNJJ2nuCrUDz0ojAXvWmwbKoZ5Mf0fnElff5SErEfGuqPlhuPEzPorgV8OLDF
pdHRiTTIBHrvE6hT8Es7JW26O1bwMB1WXx3lgpdvzh3R8WhUeWcDZ0k5dj+sEaVYNbH/O9nLb2lG
z8tP29P5g7quPXRSCGyzLhRWzZjyL4OIvIh9uouqMBB7dqiMfv7QZ6g5dhTntxNI5NaEPjuqOvwx
I6pc6y/yyFIiKeGpbeWlmsR9j9iI8Zd/XV5+9nlYxSUYawV85iqMIIOGqPlJd4gUIbWgPoYtHrNU
knE66TSCm5hRwFbhPCm/uW4rlp3VWtTw7HEisosXijkBhfduVkyCv0Y7DejEq5Jb/qFPoHnBGOK6
rOOoA6A3g+96DGpsyIxCPEodsI0YoByTNCJHUykHX4QQetlUm3Nmn4K9tu0rHY/cjdsEzpk7laJn
FwUyBrgO85uIcatJXj74zih2qYF271hzD8KNBgfLMlid1e3G01skDXcI5egUZtuWMCBuNxd7Q2AR
xPSnOCheEQPjzfyKqYm38uBznLbVDGw79xS0DrjmFV6LAGj0+Ezq4rvebcPyFsGiK7RZgiTTprdn
MelQhveG2kV5fj3hg4P489CPpJtIhf+oqKkZs1hRC55l9QOEQtPb5tw832PW+HUjJ4q5JjcOo/s0
9WnS1zGsSwMtykJ5prn+l0E8Qzq8iTfmfuSlZFQ3OqSI86cO77RNgRzTxyKNkej1WFt2kpaJt4PV
el4E0U3aweMLAufYQaCxRwOaBhV0QxM2VMnRotQuzMn+iHkuWaY79GdGbSdTednd8iApP5Abn5ZN
pH8JNrC3ZzSSomVdXJNHBUe/CxtZfgLj0YosVtsYODv8KaWhDD9KbmUB3OlioMyFJbSjilqeoqZ6
DITwYPj8KtDyjJSfVWTTAUq/JH6hUKk8mRGfbg9K6q4QfpB0LcjTEHBSj23ZkFfjRJZQ381gcOi7
t28IUc9RepAP5xIJ7dDZq831Q9WJx0UexsKrKGW59WzyikLNUOYPet3URWE/VVQYJoLxnYGZCZ2Y
Aggqj+3zAZkAvtXypYUAGPyP0jnSBJOEsudgeKVxUWo3wT6RZ9WE3DmaHqC0TBOruKkv83dV2kS7
TOCAMGcjnJBM1gNbXxJTJsoviIJ0Wm13OHm3M+gfx2/glga5nWy7SBh+11Y/JBRrs1WOW9UOmA6T
ij0svg08EKvUCVpP6rR0jAXX8BOU5wNllTza16P7Fv0wJAS9R/oLvnn0gWYMq4/wrtIyROd2wHsn
4R6EUCGXm4/oJZh4EuJcsBeEHEr/1+b9gJi0cvcp/wO6eNF7Ro82ZoLQIasjiYt7Wyi4PpsAbLwf
acsBYIJscqR0VFLWuEAnL+NDQ85v8LHcPd0L8WY4il/snNahmrUyF8cPW5kq6/M5zVzkFnbvsc/w
GFg5DUYQQCJH9dadRO6WGkoNRKe3GNMEyoP/m4oaxiJylDypygP4HAZQEh12rrQxnCcZeEiArBos
HNomTwR4tvc6lLZ4Z72vF8jX5ZObLRv4lWB5/fFZ36jZM89Jr8vVcdENd114OzD6c3l/7N/MfjfM
BD4UNBJQUMyGriEgFRkV3NSObl3dbNr2RetG5UoHS0b4llt0Syk9ay7J7gWJyGUThAVdLai2HcVS
ZW2CzRGDmioo5DNWeSGspLwNmlWo/5oSnS9mhBTVNaZcOusO4OVshs4ozWvE2RaUadDtxbaReZaj
fM4k2E5vqoEyqKtwzZPm3Cu5T9CZ61bpjCl9twlcAlL8K4TYgrc/my7lNyxFm+DYI798BENiwDwf
LXriA35Ka0/g8dxi0E2UVni/Zq36v0A7HC4sH4BG8N++GAi6cu8xHk+FqaFUKYISOtp38uWbb+VY
aQjArlwBg/PslAyeHi2l9dSBR/eyxCSlUlQW1+pPe2VVULk6fkrK4z3ugP5SVxp6QDHh9iUtZ8Xc
3eYXYYkvaj1raICwsaz3qojbmgDQWSUClIG8wY4UaJh+0yZAWLINu3/96zfWg0MkpCCOx8jc+5Fl
Q9gjAMPXyay9XODwtoNzamVyUH3Aoeg+HE7N9/qrC03FpsgIHrHDQuCsq8tHZj7OgB7GEjOzOVbj
gwZWTKpzYTg4+PHef1kMTwQOHAV6gdXsjdkFo1UKkNDTu6cRddU3WK2fRG+KE0xOOd035xhUXCX6
DtPm6uQW+8I4Ua55CN6Oyce+2F0Mh4ZQykfwS25/UpzE8PsniUbkAX4Fo+bZhpphMeosGQDPYAOI
KpQ6Tq/GLa4R7ie39zFYJsHjjVzWPc5JfdLU8g5ktBIv/yZgfMZwOZ5MSWRHsFHI/wUBvkXN2ayS
QWcy9ybeR9xLd6OasAWWY/6paciuK67FGhWC6uPuckpx2lZmbTdcxymCKjcf2JcIxp6gmXdfs2oK
JsDeHEwZ/KPgew7m/yY+O6xHsXKWemdWhsk8NriTzcrWHMJRKFGQUE28Dt7UzUKK/oHnbRDGHbxU
oe5HxJG07USe1uadz1uK75XLv8Liz0dANgGNNNUx1Pf/XL4tNnG8kfh4w6s7Mgav/wbzPIISP8p/
ZzA+eHpesn0ClNLBVJ4wYdoz9A/t118dtIwCnzr/tPkczjesvEs6phlNySEwd7TxLtAjkr9m3xuU
eMpcHiJk0lXAq3QNmS90+pT7Hlo5UcteB7iEXDIMHTF4x1SWLmeKZZTMw2h8OED39wBtWrDZK2wp
plfnS1f4/z6RY2ohOBUfc5vPUJ7D54XlZm/DvoeCeI7NBWrv9SweGprtOEEslN4/5TOABjRP3ZhH
OSOpVtQXMso70Xq2frCBWqtpHhwX7mMyFcnVDverO5Yc6P6Asd6Jc22zUtpb6qCK7gaQ2x08K3j4
JmMd0+M0Y64MUWetN617e/7VkPgKTLHykiqZOcl5HOBpHu+Pfj15pDo0Ud3PK0DvNc/STQVNgUWR
r13pyJzZO7RrHfiOHGipiGhAazm1hoMc13GolUtnp99dFAPJSc58B/RG9ugQ6URHvZKdem+5RZW1
dQpVKtT36fqtKXASY0q8N456zrQGQHI+b6zuNbzS7oLOV/lQGLDnZJvaMydez+s+QT3Mr6pRgIEM
YwOME9tB4c+VIZErPUux3n9z7KSdrlGcr0ZaVEpgrx3c1pbX2yZ/TLW5E0EOJTO3NFYcQwppEx9f
hccWXINkOgwgYW5f7KHbW5/FhHFFaRNvnUCGTRQHyWgqX0rDZZYh7AfjfEmTmY6JscTJgnMrhhvA
QQUvW7Mr9y+RJp/GpRrm+HS1aNp4sTqqE1miWac1j5lSPX8kxMwnIpIocf9QNt2xCPL20jSOR6tK
cJce6g7WqVDg457Q9aqT5fazYxEz5YX13bsQ5Ae6ndDbycPEp00EfcZz6CV+yjwqBGvPTvbQqQhy
eNi7UGRXPayYp8TbtMFEIu2V4UFI89RP1CS7tGu/sDHW9KUutV2Li/3rs1ppAY4DjtSfgUcWAfpp
Oib2czvXXeAS5nme6l81fLP/6PNYbUl452G7+XfjTa/CW75cS9L/CSCfCP8Npdz6aAq+6xLQ5bje
g3cL6pLOvjX16OeUW1qAXsuoYC4ydH/oaNAiy9QY7GRL+TnfNfIuU6llXcGWOoIdZ/WG8yaJi13d
5b4zP2HLhFUF7l3s53fP7ZJss/rOcJQuYTXXflgV5hpOZIErUuSeyxuE9xbPvhaHelZQ4A7LNdCN
EXzFslB7LFwtzPEuAhXswVx0W8ZoZYb+W5HbBrFYz/J+62JW4f2ChNSqCigqJQh9uwR35XvkfQg9
VjawYlHr0srTnPiEUmy0vU5mJHyOFunlFaYBIazaJNf9nqeTZiZM+rDbWMJhq25QIyY4WcW8b/0r
WUBPVg656xiHHeRk+chEH0B0knj+2BawjOJVWHeqcmLUzxMll1b89bJA2Tb52YGk93tpEB68GFrj
cV5YPyqPVxVqg77hkt24SP4+0zxJNsFoAuzsacjar4J5ZqEgVv43gq4GNybZ2a6hOuMEmFrTNtjw
5HgorhSWOwJUGVmRX3wcy021bU1UdoYtEXFr9dA3yhAnkmPuoVG5IR8oFybmpC25uL02seXaAaH6
f1e3sQl3pcPUizncam07HlpPV3hUwoesUT9mvwrY72Bq1OOww4shhDUSpfxT4VDfr69WdvzTAGLf
Y3BmbHr1UezHdNZUGPO0epr1CgmskUXVurKoApqwPQF/XyoWetrYDD7BeymjnrpmlChYmCwGJWLT
XSxHzfte6rVPFRXliZiszXTivhrnAWx9A8j72G0MWsmHksvCUmAOSZx3f0r/+Wap550VZEoE40iE
qQHE7pDSJtmmhKPvAQtodMzPxvu252MyiBBAhPHGGJgJI3JvR2cQFfOjGMNPNowRxXw9zdbGLyca
rGqEqtfPyykDrRr2pCq+5SHUz3XY5pAxMJCucsgDqPbcKpP0whW+WeL1t42WJHAKDsv0X4KQC+YN
tyCJHj59aym3SUPGMlXYNkPwWvgqYlmNzxNPiAcho9oY3Gnzx0J9Z+S/QTzTs22HvT6i8F+qTQdI
9OQ/8Ov2wuob6WG9RNA/F3uwmaF9+ct0HGLkPdklRDLGpkrqBUUp1hisu6YQULuCZbMfTzBjkXan
Rm2zPCLHj64hHiypp6/UXWnNKflj0uUU4b9Y+TFY7TNIjwvPON1m3rOWOmwrwAbreIr/5f49hJf4
7jT/qgWUMmoiNh8tDFN1K9ygPGzxHokAYb4Tdr/JYChvR2efvMDWjMplacAjMiie2QZBUncQ5VDN
V696k04aF9zh+Eb0O5JA3Qj1kb+LCXaexmKBy0exAezWTiX/ITb6o5Q85v8zQukhT71ibG3nfv7R
6z7dJ+FyniiO708GLt6+hCiSvgBrxVSojpgwOGjQUo7kWTkzKCEeEkHNDBVO6+LoNb9mbig7dV7D
qchYEx6ootzKWgBaJTGDqrow6fWwnOF6dkYJb5aTFQlIh2A8M5Nntw5gd+7oI7v1lyqhmsIc81ih
7G5itTyEgynp0KlIwrONtpfdBBnKhU8EdjApvYqoC5JBQ2wJngc2jc7EBSBh/PbXgBZIA5p9ciVz
kDTpEe3L9sifG7xJM5tEtW0CFXK6O0awymIY5f/zAkW6oPmMRyr4SQWCP16KbhZNk9zm77grkboD
uzbl2EP2DePTjWUBYXtnQVr33bY5kTujDCBvVqGxUIcMh/rOBSI4a3l8s9Zb+16uZF+bxKp+C1Xd
OQVPjDOhdXt6PqROKZiUQjMd5S1pS20fbfumgnBez4+BjL7BgIStCcCehd66r6c9AQZmt1Md+nTT
5Gb8kjrGXoGSdgYf+s640OIkBynZI58PjBOlRoYmJBHDTvJI5455NtvHpXaN8iMcgOLbB9O1gSJf
HSdG0vKxHmoA40EjIsOr3qR7JFqOX58aw9GS+n81V5GlTp45EeIjip6fc03hIVFgtUk/VTfNlxAZ
TbPfJYwS/ttgF7wTuJrzbL04te5YmmXQoVQQFdh55UO9mLDpG0El1pJ5JVO80QvPZaGxXJ0oNvOH
+9HlBNrrfK3Lh5POUeJgdWEY6IF8ES8rYZrCpsJhJ9D4GS7imlgyvNIwUMDJq7UtG4c3zma6TUIE
iFiQXpJWE46cJmu/kG61aFfLkQzpudylT4CFaq0Oi85IplsG8IxVVrVrOhjBKJ3PUsjCZgRpgEiY
qkgXh5ZK83OOYIzPUGOjQKU9klB+h8zoDnbruBQ9eGYdigL02mx51hGINBd6TsP+waf48E1cbIw7
KffGqpH+HW+6vPY7euG+qMPgclxNf3eJL+EoOQB57kyo7dMz09WipsEXMx4ma6Vzp9hlgNnIAZ55
35kE8WrusfXAetR0ryPKY+4mDWonyb3ClQ7D8w1mq3lFjEAHT2dFJZataHxlCaq2brSywNelsJCI
bzpUNITZbVdt2bf96GBpksvt3nG7u8QdlawgSyfxclXEB2ovS+2nxjD0BktWbo6fQ3ev6btZpkEs
hB37SCMjDYHGLMFXJGBkdUQJ9JJkTGSy6SircA0VzsEfwZZ0at5kznKr674p+AqoqD214sIU17Se
HnlQtfmv/B9JU+6iIFjaGnpopwhXggv2VU8UvoSWy3SY3SaEjx0GEbSSuB5mTtTEFRotEgF9ATyr
YVfIYrlBzvyM3R7I4V2u5JPy/BCXKBD2Glcu2FVdrk3JTeThA5pL9I7VALAro3QEv5o2N5I/K8jh
SNJEBVwn+imuzn4AkWbih/8akuzIBOBqUS1DMm8wH2lzI7BWNUrbhJPNlVtZkLnuNwiQFh7Fs/rr
2meWNTRyC/XLwC9P+oElnmb2Lq2YI95cbtLqZoEVwBw5tIVAGLYYXnb8QoUWJBj9iYs8TDt+bYk1
IlTlq6tuvKzmxzfXW1DW1KMiT6FntW4m5Z87gSOrMrx8oHTODV8idquKmVkml3+98O0kztjow4o4
QtvTr1lk2OFq8jmbGASVxpaQKMa8SXU48gfOfODsgDukXgZBvFibCquUgbq8pq+Is71RbX1sJbt5
RfLfh0TfFhFrXT3rDhsaCEP5XrAiD2XwMQz4gHT8kEetz9r/LotEub1PkrK0kxMK2NeTIeyPTmLr
e7gjS6NMNNLK1qlIQYPpupo06H5ZM2QWS7W716tWh5fatcGqUmYpglGZSFdDN0Ake1tTLr6baCvT
rTy0XirrQGmO3E7P+vmetmOKG9+utK2jL54LanbRXfJs2czPaSGloiquwfALhLB0HFUUf6EJhbsM
WCzSfhCfrLhJgUWhDk9S+QIOdxonNTIcxPPXt6BhAKNuPMxuxLlmAPSsKPaJxHHy/kGzgtvR6yFd
2ClXc7A11kJIWxppKoJGoguEh/Dr76o7eUecgZ6UK2M+/9hjs3LoIHs8Ii7Ec95IDRo6UwsJfxbp
D/EeEJ7lDnYcBn60MmkI8slGoSTfh2I7KjlMY/8rlaV+GVgqct5aOutxpQ15fmjBx0i3Kf+eXUE3
IKJ7DrTZdjPyObOGxXm4Not2y67mjaGDOWxoICuzYmj9CqK2qGEHX6abMfzhPzDGw4JNPOvAjQ3X
EA313qZRTr2rbo2DqWcql7NAsy4aaxyhqhZnqfgv87NbtP3l8YQtwIRSsQDu/LCTmWxZKh+BH8NJ
6oaSRG8+SxA4FaN7F29EzLqQmTHbuXPLkkq+RHOqWweF9m4yUeALx1Acs1TWgILMIaULjxoLzd2W
msdUAXI7WUZwysftWHJTx6yQBP/1HTgnEtpVtU7KyJM0n2iIyEjFQTN/oFNrd+ci9tgd6h5PlCNr
02scgqUZodkiNBdjeyYgADTpsVMIxaJYab+iXy+T2IoA4jpIrl+flyXSLgOBBoElQWplCIZ3IIGh
v6g5Q2mQS6jVsPUTPZ6SV0Vt4iCYziSX8+kZ5JnAE3wok4/YDiZ+srtCl+RwFeyotraG4DalIDlw
8YITiIwDrORB/aokl2KLHUfIgOYdvL8Dj3MswfE3SPwBCTScCYl5QjaZc9axE2yIqb2vgPPdU39u
Ox90SeOgM6il+X4Nnsa2Q/VqKbV37kLqfXPUdKwJ2+MsyT37Z1K+oMOqEtzQKAe8P6bNgxpUDunH
vcZiPbkaUBHHZQFvbAfeGUwUgiwUg1N1o/D0P+DxjBo8Q7htzTWp4jIKdhY5vWAgVlI4/g5jWopl
i2AFyfL2VFo4s1lAYuG0UOFMWakr9M4onaNO6TUGDDCrx6Dy+hgQsrNqIstZEkGWEnAPCGxT1OEX
mBirpGxdKIMOVbtqC9S1gr64H6TCHLKUTs+zfk5p3fUwik8nERQVPbnBCj+mMRk/RwEy0Prhawba
tUXBf+mRtmJzn1TGia8R50hc7NHfirgTiSHAdizDXzsZvmPvl1v+dTJ3UClij1eKF6Le2Z8yCN/c
MQ3s//zrLd8A4bUTgGIIyK2zxrFTgtWWIvvvR8H1YKW6GQVF13g+b5NafccDHP02MQLPRoMx3NfE
aF5Ww+rl6brDvhnPQ+5Q0QJf5I4QRqFQNKpGuqbBVeFGKoIPVaJauu2/IWyx1EeCY/zpVBIt5c5q
3slBjozmHuFPCLZKcUKwM7bD9DU6YRO0ubO1gHhrXT0TarciWNdC/EkI3TURPtg4TaF7L2o/VWxb
YLz7GEhsLFloIcWZiadE+1DIoUv4vlVbmQ7RNATAhVreOl+gDPOdVRxJm9+x1GGTuVE6k3fysUY4
iQvowdOSK9ejDwaggWe4niI7NcEh1guHzZsXb02zwUvGDFGfTbQOrFTL41N0AEv6GvygOGSSc3TA
BCfU39D2UlYekjOXiPGZkri66sMrfbLiSmj1u9UYV6oj03V615ihz6f0LHYfa9oyC2UBox8Cf88s
/463vB6Vy2CqUTTe1BXRduFd8Om75rG0jmXixiMZkuc8sQJkc0o6uXaHLMxZWjXAeoHd44KCsCju
omcpOnPD9vsNALpvvM9DvZjT/Zz6tuNaWq2FyIX05I4vIaIKvR8Q5uJNxMPfdVy890RHKSu4Gad5
wIrT1yG5BbhlWG+5PBVVk2XMOtDCktw/avtZ/upnrZzBvqcMyC1oFLp0G0dCIszrLxouPBr+W8Xv
CyT/jjym7zwijK8G+q0rcnW1oxZRwzKjxab2WI/7BsJ3OjNcZ/rp5tne2fM4SP0lLg+X12HdS0+l
1G/r8gX9mo4vn4KiEWDzGrT3zAx1/Ds+Ck/ZA+RM+aEkcynL6t8II+spXF+jzJCOWeHpk4ofxSRC
IC6wLineGvkGugtJ3+yG+CE8zbr3wnA9jSsfCng0QmFfwGyJRykZlPvAuTJWJmaEyDWPyKl/7x25
qRa92h1gv/L74+EgpWbuxTtoPohR42qiByXFACa/z3OcjuNTzZ6Ki3o5uJsm4ZpYlaY6BH2+JRnp
840/X/UtphNMfaKdk/Fw3k7gGE4YBrOZbbq4haGacw5jUJ7NhSf9slI+zAN2VG+N0oL8/yojW+Gu
gkU2FcHVlAkUr2yamiKviDm6vjYWIy5uEOtH5u0gphPJASAP6AofFcd4AF9on4+84m+3jwJ0lLW5
KcnXqbZvTRtWCg9vOPvqOCcrFWHDgb+CH01PP3uo63Do9rcEO6gVKhlSRW5CMkP/WJczmT6sMApP
91IXfaz+QoFyrQ3KoRpb+91ADYxFptCU5qk26+siaETgGCXRJtbke+YZBEXAsQ6RTQr6fR/ZQKCB
ITM80z9QRThHL1HnjZyRHuhFbUOYIDUf17uyx8Et8S+tfGQfNBayafSoMoS6tAQlcFSmW6CAbX0H
ERASh1iOF/0v/lgHGdZB6FNv6guTTPCx3TuyOPb0uVLxc5Vbt2dc8BEXdWBuyAs2tgawuZNj0jPS
rL45bWgxueScQTxm9awSDYlZ2AWwKY8qioZth+PQhEVfIaQlUgQF10FR81seICT+QiFClH/0khsQ
zgMCEA6T8pDQj9eOavfcaHaFqY9nI0rVkl2KRIc/oemNK9NthJmu3x0G7ZNO8vsxEMMhIi/zz+hi
72JQfvop0fSfziHLJbVuXWSwo4IwJS8B6LXS14PgVPiWrx7AV+kF8/WrZiXsbgzkMqP1RArYIiD6
Ks7vj2OI2lveS0fN3KdGCmorbEmv8nWHAOTLICUcYSRolzDfJMOOrwriEeI4OZlcXXYkqnoi1Hio
wmlWcMvPAPlndUuvzROiAngW1J4TFNAYr6m1L/1GG/yhH2lRm2P5ngu6wugypqOH6ivK2CWsK6U3
mOU8AYvlPQy0THhb7rPCK4oQxFPYOotV8QNZ8OcIS01EnVSRA/prI7GDKdHFDgcHsshDMPF27H1T
jzdHjRVIw+j8Zkffkx27g/xUrc+DIxbogtduuZ8Dd2+HR+rpYtd4Dx+VBJ3yWyDOyJyt5cGlKZHx
uycxNiOBp+E2ciOUPXNusQkbnPxSp30INMwOgG2fxB9kNHbuudsTHjw6vyywlyMhFaAH9uzQ3cyV
SsPYVA6HnaeURd4vo0HRjRjoHCdmIZQluou+ZEbuFOk/wfsHJkg2V89wzOQHD7DOIfJgpURiohzN
cCERD/f73AofvGNOhBrK0Cbq/dn2ivd4AKxVMopGvB9JF+S3OyiI2R7daCN7zTxyVv4kh8oBtTjW
or2ZQqBi2xRiLi7hnB/fEixK5tZ++T/Ei3qu/wYpw6Nm3ESfEIx7iEYx+HyKfztkpFxweCjMWzfu
W80v8NGVURNMQSJX/kdTeBjCxWE0FoSVAoTKJZxmL2xaoHo7lCq7E4JKzuou/Cej9yXb8qvONgZC
QU7v1TdNpbFpdszyCOn5SPHWlrB9jNRiovKid3+MCARnAV1/zqypSrnXJOfIvRKj6LnCpAmspdV4
S5kRuAsHGuuuCj/lH6GRka+DfxQEcaltxZScZY8H4UlUt2YIIu00iXny2bjqfvSmHIaRktCktNN4
GJ0LkbbyEykiSu19re2Jj2N0VtxClotur/E/OjggcMCxJU0cWudYIMQeU7FgxpGMxWAtDi0TlRLf
9Zd4c1R4K0GRjIXHsgmiXqmzU0wWQyXSo1rZIlXTER7Gl4fqZYn6t4BhHR2apflH6eatd5/x+Apb
qx8OjRYqAjo7C90gEtK4LqA/3yuMCdX89mBCClTe2HQBrSCNR70NTLuSSMAIZjmN0V6xfeM8R6mx
bvIHcHCnfKIsGfg+/dBWdeifEwej4bnd9wUs1FFA3osajj5VqMmU3KBw6XaRd7+z+Z0RCVAPYbTJ
z+qwh89gvWieS8bgFz6rnNIDLfnE4oAPpuj1NRb8E1lT5AriDM9ybz+WXbCJ1n8VGo15v1s672Cn
5VKD11KSPfaJvdPCyzOvZBnehNP5c+gaEQb/DTjFHt8CH2TKxzrmXqABk1VBIppd1s8x6t6HHejq
M1hPnhhEeoLs640NdhDt9hvzGKHtgpROHJAbNRHb+6emvz62uVjsUzztqooZ3da5yBl/n0MrpUdw
PuksUi244WF8zTBDjrV5dskZkIXO16Yw9VPRXcRaD6d5tX2bFCP3VzKpx6C0A1RxWwUcGeoPbxeK
fgJFv2JClRaMsR9SLTNddZqWKcO+pdLqc4dHxp10OE5j77Rir2CXb8xWSUqyKI6Jzv8s0qJWxDt7
hayrZBiRZ3VQNgsBoSXA4ZxsjkW5Hee1lvBmdQ60KYrZ8dYdWRmBtJZMw5I6fM4I6+lY7M9G+iTL
q7qhHqYlBurFg0vITJDx8A8G8sZf3K0b7iy84SNFHRKnJxylq+DEDn31RTgkS5hGIQUanjXfyi5l
WiefHul7ICiVGhCtoi7dPlmR/SHGbza7B8NI4bqIMSG708Q202hfb4IG5+tF9YepljRFj3hV2ChJ
QxSSOQJ8aaa6K9BBX2BfuW+vqKaslfRa+I1PSmK8w536lba228+Jl2hpbD3nbdDnmzyti6FyguAs
D7na2s2c7TG1NffP3G7HTZPvZlnLluufCo79+QqvPcMTP7rN2oX7bY9ElxWLvJDjYcsMGo4u/kgX
V8vFTZWKwzBVEzk3+1w8XbwnG7W5PU9De/CXQXdv4ma21hYqukdjQoonqecssyNt7aUk7ej37OaO
wGKiJEBtAeljI92xWHOlSkFc2mTepSUdNZwCf6ZpYrjiERPKqTNMGL2ext/w9cnr+LyLBuMIdVEv
F2/QpwNXWG1l0HeaGEy/Fm3peBUVWOV7HnDRccBcD1jUBTZW1jfN76KUA+eZS1sxW6xck328DcZa
XQfS91+nyOxBFXBoa+fJy6vci97LgkQ+sDn5H2CPYhntbk1jwGz6dMERZ4PiFHLt4gjXzbUjAIIM
GW1jmGrGL/zEC0ucGFMdwY03DGa7emNAsyrbev+t1aI8neL3wHKdk8OXMhLUVYCjMPaOinVQLLn5
Xqyx+X/bGQRdqHshArL4cHzexd5YRB+a9xyIi0D/Ju1zNQLNyCRIQBZo4fXfbzGaGf+ZGEx/FHMF
y8gx9QZr5I9jJmgiTdO0ASiGyOJW6YHHfDodacocnhDWMfaaA/+C7LAGEOxZb0ele35qjN1Aha0Y
61bytGQmgN9uN0VdP3PJu9ToyD1tCCoWcw8Jq7tyMLCYuKsEGsOYdU+0XEm6cJykjJ6p0Uw6RkPw
fa3NxEP0Z0AqTjAOn2EcQlTPeB4NwivIYGmvGB5OP5enJboCgv1U/ug79Nrp1pyM1oVzSaWV6NvV
2TNywiiDn/q9FVgqB53HAwKvSyZph+wJnehKfkEyE8FeA6P0jg9H9ndZlEgTqvHQDBgnW0Fosb5q
ruj+h7HpK91tilmLS0BKM6yomcXmLt9Pmo22XCFhzoIsw5zHRAHAiWmtrhuG+5Hv+6NJgEYnR9Hm
zkefR9k+HJk9V3wHIuhFA3zcdYt12QAUeO20u/8vBWkjj/QziV+KY9HFqwNp54YCv0b6rDx1Rp77
kOVnUjBiwbTwCMVbq0XM+PGtrbSJFDwuHH39tuAr38fkJCNLC3KDoAOFd7FwI8k3LKaKN5YnL3qZ
25rGRJR12KAoek/TJYsdSPeRP1x0eTmEOcbf7LvV6dOKOtMEJnzA3OKc/jpcZSPRXgS3yuMqLKsX
XeKIbURb1WlH3aD+px4YWO27+FJJRiShaqnZdC0QUce42m7Ra9g/Zs19rkKfecUejj69wZP84tke
ZhFm5LPzg4HgJ8JA+2KGlpnV3b/6YnCrts/c2PmjQNmrW5No3lQrmbxqvat93XYbBYy/CIhOBu74
h/e8T0/NLhCe2H0zdyEcECBLgMZhgGINo31nO74+Da3rTXmx6z9V/YNBR+EsYeaNZIBdCZcQyW1h
mGuR18zTMRH+fKq3fpIkOyTyUE159h81pdQohrKGO7PMoIrGj7t1iY/vAXF8YpYpL6LZxcJ5hnyd
SK+3k3bBJXfC4+WccQ1Rv7vyBspRuz050WFbu6WNQuU3x5itdLW6JHuixmPJeh7HIXVWExQmdcQg
26P2s+YCTWEGq6sAu1HuYXj2mAl98aj1CRBBV3NjcTlDEtt6hEqjnXRISGO/Vj5Us+XYXeTEVP0B
voHKz6Qh8qU+d+Zf7skqsyKLeoyJkvlqoe92iADDIDOuGfNrPxwdYxVZumGXHRNKKKsNzImSV89f
6vzBJnensLqZV6RLzbe0bPNkNIQJLiUwwp8jQcJ1AIUPybdDAyh4ztIEKnhTd9vAXkZeM6sbUe8Y
4LlP/x0rZFfB05V0KKlhxyM467Ia/EPcOQ2e+WOWwKO+0zU2K7k2fffG0mETyykfoIdKkC0Piwru
MwwBRGes/HvFb0Z43sn9HpwR+P+371dS3iatJGxalxptwLxKveWFVaw2Dj53YgTz+zJiCBF7hZG4
LKZ+9pl6C/fmNvJJ0hqH1LN0U0Mlmo8uavWAEcDB1Ocj61JMSlqBk+P1T+XoYKDnKwo5XGWEI9eq
NX44U43D9R1XEXK/apIFMeJkPdAd8zQbhoV5h8JAqwIB/v/1qdC78ILFJi+3Bu6T7lwBy65B6bom
VeIwDv2rs3W0X5Peon7oCSV6V0rIYZVeW0dhlV/JBpLn7K26KBXdnLdzNdIz7w5gLLulLdFRdEu4
yVWOBEdXSIyNgetQ8xZnSd/7mlEzxpjhzZwjPuj4aGC4J48Lw/2BJW7ZkfyUetK9X3vrFrLrVSB3
Za2yc2oAZyv3AtPR6b9nfFTjQwjlpaqI6Z3jyh24jRqo/L+aSpQqTjS1MIGJnE2s4s0aMp0xsv56
wNgYLo9e+xLsD4HFLK+yMisolPQSgTCooS1TmXDOQ+DC139bWjOmwATg8hiz3c3kaXKIrc6YOxq/
SfOKdndVCMklpcqcOvr46DCURj5InkUCh6/3BOeLKbgNXGwds4PydsGCEBX4AY73UpyKRBrNp9lG
ow6QYjw3wK+6ruxH6LudRjVjB6NYdH//eLdq6qfAkqLsnBtpovxL1LSiZy/D1kihOgHv9aRqyNtD
Fn46I4XZ6b6+pKWTZ6y97ddW7mLtdW0+gvRcluHyN1LrruXyI1GMiTMl48OLv5T5S9hjaTyMjzj9
TGYGcWez8h+THFA5JmqlZXyHKYZ9G5LoxG//tRWBk3hIOvew8nFs1CvgEkVav970Z9IUD0W6Bsoe
q2pMyrvKIdDD462+X9jOgP0x8tLA+FSejBCwKazd979nvfIxnbJwEJUDBjpVXu5ZcqQkhJ5mYnBv
KNvZbZh5mQjK1gkOIrQ3t6DSqAWexeVajUyYJ+tjYYPu//UROmukRbWOPQhpcAp7wpVhaX+pVE4j
/myo2CImu6J5cVS87ywsi+u2kbsSRFs677qCVRkkRekSDSJd0yADXLTASjcNSWn8U8E6iUmw63jO
GqDj2DJH2gOpzUc+Ajhg15VUXOyuss2Qx9DVlvxOW6Otlm3gYSZZpfUDzYcP8fKtpwqGMWUfQCGj
uIP0dRSIxox0sGHK0xh3s4jYFPRGpj6ZyJ9O0bUB0eCMcUCiKqi0F7TE5hYxjJdGeDifUMPCxpBr
yem8fjfUmDPwIaDe7+fwlcQeCVu/lXBxfg0eTPFiy0yUolDaIK4W64rXpspKFTBCaW2QhVAWAvX0
SfGAljC30J5ncUYmqzT+wGB9MtWtJhbUG6k5GKU20Lyo41Yh1IJYo+EMpIcyj6l7Mrr/dKpRdqPS
xD3OPvoTs7bfw1LQh4VF+i1irRKzB34MQuXhmMkMi/6x/96BZMC31jdwGYGaepIUsKqM4AUhjjTB
YhjuAL7Sbw528bX4gCbBZEUM1+RJwnVBt6apPv8xlNtJPxDkyqwXOmaMbyIc7iljGst/zoTVcS83
hCeZsas2lvv4FfCrLbToYFo3BI3j3IGjguf8TnvGRUbVpZeHFztFs0FImN0LT6IkixnJxQEKnGVP
PBVVY2PYpD6oVrpw/YItqwibUVdC7hq9JdiOJwXG7D1B/CvkbUvkDKR5L7QggTzu7CBHRu0J36AW
ad+i0O1LMMSVCTQVjrR+EZK3XBHp6idk3rI3VXfHJZ+r77/ZsulkHBf35nqNAeME+rGriR6k+s6I
WofG3OaTgeNYp8IDGfdSmwl9o9xpA98C01frUCCYf80eJHHdExuusQexChiOfIxHO3XRO0mHiFtn
jwCkdo+G8BwTPvV4SOSqKvchY83xgOwBLgltKH4TA8AIBZVzsmPmfOiKEVVuBm6CSxNmmUR+63De
EqEueAqHD1I7bgbRUwaG+OZ+yfJI8pBi1U2upzF3pZhjqxrkMAvyLH51YbYUmd6cUR3rbaO17I8e
iVaRosb/wQ5cVRdk2zzAKP1q0zQRI/pFqzIJkMN25h+ZrjC0UlWb0vZFEAdQ54IE5nRbKb4wskFY
UZAu5TwPX91MdvRv85vlA67m3TP+1WHsjN/pUcN08ZpxoWMVkXQZQxgH5Zu16/15eDEnzqcl8gDQ
OulfMwmLhd+LSBHD7VwWbaOwqo5mBiY2kJLVKfkpnPxLkfqu5PPx/pPVEqD1dlhXPjAIgMonkXUr
kz/4FzhKjjAzGrSsv4pltMlnYzkU7EoiO+fsj3t/BToP7/zszhacgZK7LWtC1sWBjUbFnZVMhWvH
f9NGsm2j86uXqPqu1AIwvuEeWf0RRH/IWUJ9wZOMipWsqAc0RiT4IsaiIG9d86hEvKYOW6ne/y84
+Rs4eE/6rb9f7Hj2yWDu4h6VHPFbMWvX0Hu45dJJSMpoPT65aj4pFtsFNV1mSaecRCrxtEvXDy1O
Hhocdg0OZI41xftBCDjnGg/Qx4lpmtsZgvjQDFZHqO+ZFqvBbqof8UV2a4UVCMVJRuJS60THviXI
N64sBkwBVlWbEnHPgzZgJv68QPAw5A+/GSGwZj09PY37W/nStB3M5qQd0Gmk6BMyMzMd8/Bu/s2H
bL33x1RUiQi8NQnrXaqhtaIZ/wXveQbgJR+kN41/r9nA7KC4Kd7VQtd0GgTORT9ZUO3goKgYsRtF
BXPIt3Rdyj04jco0JOvcNOscFqOq2LJK9/1QckBRAY/09EN2QowJs6Zwu8pxAXoGEm7sqE28nwz9
raQi+qBEzFK39RwbeV5Wrll0xQWPVUjhjTMat5W7xGsGkx9Jn2uJ9oJS9U1dKg71mhnTVfBp2Uh1
r1lgpEnIcTqBVuOsK/pNpIiGKuhZyc6Yc50qXJpgJtBEcxOGQAeInzKwO1hpQXMijALoXHByWKXN
9c3Ek5kA1lLzLRVI5+Ds7tiGHQWRCVq58IwG+wEak2p8qXRazEVN9848r2ZQIn5XS6ZxoOTbnR5E
nSpq4s/HQjIVyU1CE9mBSOUFvQDUlbrk6Wgq7eaSMIZCc3LhY0iYVGPRY+oTdZmdr3uCw0ytpbgi
WuWTH1xfUSistrX+AK8dIJAzNW/pI1X+uIYPlsZNnzcRzELD2Fg3lvx7WFMh8WARiKnKhHqmQgiu
LehHyt3Nxpz8BsBE4X8fCFtBY1/urej2HgQB+naNf/lmIW7QDOByKFCYAzMznAFl5+ea1AalyDpR
sbQyJ1vvvnBnkSUcz/1rzikOp/jQ14P+gH+NsvuRpCmW0d2XV/TnBlJshYjFdXE/TyHUepZz9IUv
khLp5LpMljxQ7n462SG0jHUTXoNYng+FOE3RKxiUBgJQ934G4iLYokHaJvwrnetgsOKBshzeUlob
T1zFcVdTodv8nq3zGBbLgjqxw9tX8rdpjQh65N2IbiG9GuocKXctHEU0VjrmiMn1W6W+ZrgqWbjY
S1HBOsfRwEssPBASGNBtX4Pt1iKSLVn1Fra4nnbQ0ATyN64SXJEE4TnJ4r8hR/JtoLD2/2MIvLK/
VegN6OZQpubZTBXyY60yPgtPMED/w9MIJqumf73TaqlNG/S6RNjDr0mqoWppEUsckFowztuKQwPb
MVF31MXbRW/inUfWeh/A+GcpQzqb01MPwQaaxIEgmWCD5DrTrcbdVOz6oGIjsOXEr9/jYicQuMTl
vuSgAmCEISqxPB9n1VxOjdXB3Qa6KPqrmdu6aIAMC6qA374xVH1O3hBmC6IEw/AgEng2Sp6lutCQ
0dzap8/aUsEk8m5DoZCxmDFttSRxiC4Ob22BQ9tN7+hfEExZ7s0KFOYlbroa6RYTwtawiXVJya/U
RsH/07M1Q5kdDGNjag352I5yVJybA8OFiK5b6CqFRVlPoUnFU+5Un703XDjtDizukutLadYGgG2t
Ve5fWxqQFzbpxb0b88Iw821ANdw5C2ZtsQYm4jJxieRI3XTQurWelZrHDjMJtYTuMiuFNGezif2V
Q5X9mz6KyOtuURF4auW2T+VWl0/cTjCMX0Xst1Qooq39bX751D8V3MQGBeNylxACDBGvXs5GQ2Zt
Amau/AMY23ZUNJ/OAYAhgb4v7XPgml0ilDYLsswtkeHNGjHMdCEhZ2WgOEN0h4GPY/Rtfm+JfeHf
mGbKESohjfqKsiIn8A6xpB6h4YaGAFiTjmOP6/KIZ4ZNiNngQnnwwQKf4S8TbPtqPYyP9lmeHoT4
+QOSBoHt7DRwwKZ9Bk85q99iXHAIqdZMjA0sl8WyhCax4EqIq1gb4OWglByMrbzIkoveM1+zc0tl
ZKyEGrGxTVYUL+bHe0sA/YHMdIoYLT2lUbUdozwhuleBE0+opO6tE69pFB6Oyv1TM2ZtOzf24g75
JuBkyHi17YYMiQr1VEWEqpeh16N9I9JDV2KoS5z8YisHfDAzkdQJ+RXcO3CQGGaFHZiAvsQEEqTn
MH8E5xaqA0Uj0SfnGiIvNs/0UTPJ46hjZTlfQ2eUh526Nznn0ENDTElPSQynhTDxmv06S+EEUz9w
e2V7kcMTbNTpViGhBx9PA0SEoJ4jhS2Ctg2SdxNLIb0BDc/phaP6HdrMg2sVRFc6Ltsf0WUX96RH
ZSaZ38+6KG5AU+7//V0PT0cCzNta9shbE/LZOWaLH0PvTZ3JEwLNY4Lr+NkdtdGQS4PioS/8YOFw
sgP4j4YeC+DAwWXRykjMOoJoGMTWKiZRAP/pXuDhU6SASBYXBrqLkgMripK61pkoFyrvWN0cxAOU
pETcCytBS55pXSZPYAd/q42jTRq6bu3u6sAOB4P1QPQyPh4hFUtGeDfD3ovw0M+yZJYjawpKYbZ9
gr1k6IUA8GyYjvGngEmc9BcoZBh5hElxIGbmH433PrOrIFRnlEnr7FoT8qcznwP88pS0Ah5XMRc/
AbefSvrlOtB4jooyU6Z2lmrTSusAdvuAiJ+INXtyLCV54qkBrL2h+liUkC6rDPlyHP3ZwxIy3Qq5
RgaXXhEACwBGWbYGgMsyN8YFwKUK/6+tmg60KOF2R+l17e37jRZIy7TY9pvuQNM1OHSQeg6pbWpc
uCW2FgDsA+QJqvoR+i32VfIKqjCm9xqaaMPd55OLaoqMvcs77hrsKHoBsvzzNutOQOuAo7X+RlXw
DDGAKsjebr5qPwRreEgCTPEL2WFURt1eH10icTGkePcxrXde82AbS0eQupS8EuY3t5myI1hi++Ig
ZWedmbpync+/3IWy3TGzyyB18ztUl/+7ryilJhA0sDaH3lNBc07bJyKefzJUav3VZd5jW1Ecmlm7
CV6fRJsDRmYwoDo1UoWbYroomup5R3gTRS1lxN9c4M18kYtv6+X0jegU9cRRtwRDW161bt2dhfNj
hkUTQbadsp81L2MbmMDPtnSnaC6oyxrJ8obi9MH+Uwbriwgir8oC2vadCOS0B7syURnE4Au39m3N
Rb5kJUDRN7xH5l5GtLMpbXtvO3r1Lc+CAgj9dxnovvQ9oq0uhIe1g4b4F5lQ0k3UOfns3+hcjpFI
f2HBVE3VzQ81yfUe
`protect end_protected
