`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PIa/sTAaBgrRdRgZ/UGHuF78w31pHdD//4Ll5Ekj6Vj7XkbQaViUWuX/cqg4UHtr+KAjmOeoCz20
vJcWzSW/IA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IS6U5SxF8jk7Hz3s8j3j0NzD76vkG7LEEMqf9PNHwKZ5BGcaRwq6hAJFRJFIoC2IPq76eBdWSNMp
gZu0lQTOvXQYlsqv0WsB1t5p5uiDesPr8YjPxtd/4rtQVfHzApWRKJy89KLPsq9htd7mPbMWbzoA
fClv7FcGtDtMbH+s7fE=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BJyZoSIovIsqGHpNuAGIZ5neEDpJC/DhLUfhN/CSowWhhQDvRIdoXCnU77HyP31aneEtRsW8IlSD
JXENApSWeJ2LwkrCeXrAseclGP7NhM/xI6DDcbWxOzYZ46QapRUmLP9RICYTYhF0GP9WcQP/T9ce
5ci7vg8ujT485PaUB9Y=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VZJNzjeBsqS1FnN/zHtybYwWu6b5El2U4YhmgSoESpfH883uv30kFsDqfPDaTR9MUPp3Re6R7XeE
B/52+1IWflBPT3bCdKIpc3pqHULk3i1jvPvtXsqAWt+nCdPgyZ5eHKGcDu5EaJZ2H1vOrB/NsMK7
ije/ntoEHn04q0tieXCGeoQKfwQOkQWWSrvG0JOLRhNpr0y30cp7NTiXhplOdYve84VIL3qaAYfF
YO44LT49YFbPDyPHM3UCVTSCU8VdyFtEIKDHHNv51GUvSzK9Vw976CjIRusP9PG83mWBLkTrLZhW
sWxLFGpR9tTZIX/cFYnk4Us8GDAy1QeYO5B8Yw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XxR6c6FboNi+aJqZV2XBclrTuwMSFPAqr+SBCDz9zoxBZYK+0fIde2gqGv1kYiEeqkUvol2TlyPS
apZwLKoc/fkOcOUy6i+Oa7ektkWYibmhXnoKqtElXv1SE2DDraseWR02/bDKzBsAfmTJiTyHsx3Q
EddpwioCsJzeDfCfnAlHV/cBaiUiwYkmdSXZQH6THXFI4Xvlt1M+9JS69E0sBYZ6EzNWUNB2HqQG
kagRxKQ9uJRwTddSiftQNF1x8IPAl4/444gdVsKp7+ZLr7dznGIcd2gHg2L7mFBhQ6puMRUk/tBr
pdC5zSSZvDOTPAS1vYIFJxqC94xZ7lGmKdleaA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qQOvN8cvgpCPtPMzf5sFunRtPPPXSxdfciX4wtuzmF63oDbQLbnqYR6ym0DtlOiU5N8riX7as6vm
198yC/u2T6DVf4qVvJT4Y3uHA28LzfcGSrOqq3n09xk4QnDx/GC2yQyGkRhpVrEvU0K+IUO6fmGv
91APyu70oUm4Jc5GpMqOOusSdOKGHQ2mTedcxd4hkhmQ+4FTSdjQAbDFCSl9HNgKRJSSOq1MBWI5
K771sd2sZUCcmfFuMLjR/mgJX+WNIrcSURoMFbxJSzb/n7mlB0to1LsZBj41ZGp3AmitNj8RoCQV
NfZABIyZUEKOExb9PH9ERaWtqw2qtUMeSU2fOw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
yEdbxrHfzpn1zHakkuFyoH71QSyPs2XzDWKEWbzN2OK22GlDuO27GxLryrrhO9hndsdj7GokdzYW
M16KWYv4MIoldFPevtY3wTdiEAFRi79CupXhNye2RThyBj9197bkqBdDAD7eP17zA224ptmjY+mz
NDTWaQNV6f+aqc3LoI13XyXN2RVUcIXi1KCsCu5qaMUKUXBm05khUhL3ZBdgsMsmoNcKhkDLwf8G
kRWGmN0k2SMQM3kQNH4ownhzPS+xFHbTr9Z3ZwuVBzs3fI+HSYAEvBQ1KRpZiP2YMws84ks4eWOG
K+mYOo8RmMRRB71IWXq2T8DH+bhifrQ3rQWsSY45ri/WBGpUyvjsgw3VU9/iZHzrB5ZCpCbC1Rdh
mDWDShMXdqCVM64VGUWI/gHPzwMN5ZnJQJlrVXzEo/D/6KY7acq5iLGayJKfS7s9RCg3M47s5ObS
Ku83UjJgj1zlPZMqfkhD0fgRCpQyZ894VMcnQGkOCquiXy/Fjm8ZtTcahM6I9ifV+0pgfMLJtOCv
HADpVN8Uv1DpFqUn83XnyEvy/w0WSM/PbRqPSFAddQbhITieAv4SozQ+ETeYRaiYynm8y6PgHRbA
qCZaXYcDQRBevaau7ZqvU/rRqKMaZBFZfeD2QMgoYmKrdxxffGQZGwPGhMjKYPvzvEZLXa3+2Igo
vGJ30Q0oP9K4lqtYPODOgUE/d+fE5I3mzXHRym1U3xw1uq3l8+GyJK4MZF9vTJpvBDK4/VzPrTWO
0GCxqcqzj8bDin72iWWWo6gd+voWfnxOmBVYt3NJDYUWgSlR60vRXm21LuijyuKLnmqk+JXcJY1i
YDIyTz6YXV8+eq/Ronud0ghRN4oosghxxQEzucw3iaRk/CXu75G0NJoh0pHa1J/0jUvXh5onoTJu
UwbaxV+O1CiZw7zp7nHPUL4vQfy72nrY4BBAaomn1uAU55zCZpyfiimpOAf/mV/qGAdhLIScVi9X
qnSqOo8S2iul1b890oqpz7hAJ63PPu7nLKFRbEnsZVYDkKNiJcX1YuMPhz1qyqpjz96FkYuMEH0q
cgDIrQV1CjR95/sHNe0ebb8HLSOm1T2S1BxznpHiovEMe8x5xm1W5sNHN0z64Okz9QuAJ4iDWTBk
PdPxsO+J2+HG32F91ljPtik8CZfRjTi/fKqn456yA+wx4jO9MfxbS/CC5M736HEVsBcyoVDJfmQ9
2h+E7QTwM7b/XRLGLXheVIIA/vaRQF5MR35/hl4ORfd3FIe8wcGb8mQKSDIZxHDw0gVTYKSQ9mX8
IZFNW/JOeeg4bz0cmkHEwXIoPKIvgfkNq7up5j0486ztEuC/8eN9RKiL6s7EpLrWb+hk74G5KJSw
jfycIhpMOlxXXwWa3TEWMVXp+AJ/YSF3it85rIFI3RHNImQVcQUPmLoIR+nmqOgHSrIhboZIwnYr
IVRFBjIp78AptOfmktQvmIX5LAw0m9iiJ4P9w3N9ufMENLyGEV92cKnLAjUrI2bl01z3tWN+gS4M
CElY6JKchU2cTEQCDZEXXGxkSBJiO9J3MukWAvdTshLGkk4KqWk4913Hq+QN0G08+FnXksgKt35P
80MGYn71r8rD5qyrXEwYOqYxWPSyC/e7gMybkONnk+5NVJGdsavxYl4OM7fJS+e0tq34hVqgC7Gn
s8pIQoDbceAkXxGvx9Ehr7Jmqp72uua09T8nAWZ2JDAC8lTmNPfBZLyjaCxfupIcyzdqa9QxHhYl
l5Qtsd5P2JnunSPaKHWNvpxlcZkwX1pHRICEqNUO9dyQmPMdpFQ0HRY5Z1dX+bw/7fEawR8TSnG4
T7GTyHb7AUNrlL1A22HdV5Vhv00L7pxywnBrERNO8PdYq6JB7l4NGm1t+W+gKLTh5S3RqI2NwbxG
+qRKQ4j6+oue19nRxGbGG7vy8/xVfOUd+2EDaGChxoRKquBEQyQ5KoVoy5x5rgkV1Za+QZAruKeq
sIQkEHqbZLkgAYjFoHuHwCwyNC2BCmvd7dPwXi+8MwAfLyjrcCGdhCW/oniN35XaVHZqwqB7515g
Ce76z1yDg7RSXinFSRgFbyKrD1EdvAvX/gks48TKjs1bhNDAvJI0NFe/SSXM8L6TcnAgN4vtBpYg
uq6LQ4DqAyxKCAsUe2VKI++M+5MUIFJeihXuUjouY4+YDFerH9YZVMSUK2S0lzFdC9pndXmIpJ3B
ZFTKoivaMmfn7dsyWGzjCZt7okyZWmsLymBkXWfS8U1o8TrEW6rFTYJz7H2v85snqVPXxPgaoMTH
CMd2zgTnEDjqg1712kpKgZJPc9esve3saDFbX8mIeGOKn1WIZdcFvBqEdemKkW7Ub3WOz2jnTfte
mjrxTVHI1zE2hWHhf10hyPlD9sf5WvzBU8VOWyKDWytUfCYVbHD+JXNY5egZ/qkIN8FNUuV3nvxE
I6G7l+6rjklpyPjU1DCUo3Y5OgfKoexoD7AuFSOIpYzKwGJFhp1MX6fHIjGr4Ib7wec21vF8axm+
G2+bLXB9PmNRkw5+4ypYo7jMvAdx2AruKN/oV9IrlxRFYKM6vr2fuRiGYLRU0W6/elevtpK9agSe
7mjlKJQXt4d+Rf9mMfMEllXGsz7i+0EEpj5UX/QJn3IQWFXeQ0YM2PwvdAE85Evs952BSv4a9JMw
CykwW0MrZ8xBjgJLcbAKRFRQVLTllHINBETTrrb11dO2W9YDcu5JMwxFpiaWbUcwxYyUKjwIhCcm
QfOTIRV32AoQSVA8xV1QWcmpSFW2RoQmfAaNB3LumPxQ6R43NjbNS68WpOU6vgjiTSsNQi1LgVll
mTnvElQ7YSo4m/Q+hh1ecdPhxC9av7i/jQMu1v/yhbXQMavoVOQZ72T3cooxx34h5EKOtVpjLSjR
auvhjrzhu7hyP0tuR9Z6sIPEENsWc9NjzY7lGuOmB1ICQISaQZ7+OBkqqwSRnFEKh7l41WUtaIfM
lyt/1ztZV9qn6oj9DdbtEi2zWgnTqgPuuk85RzIRMe+6o+UmCxvu8X77IfIN99AqU/0U28i83alt
4GqBx6P6VVgdAc0UG/q2tWYC//1ebl7ACWgD4FsUYkAG6xhXGkILxspDtDPbd4Mgd3ize5JPzR8v
CY9lB6EsAjZbthonzJlJ+oLjMSXO3LcZpNQ0NzpG57WpC5rxgcOJF7hu1JMy7e9aKcJrbjTtphpF
v3FiVG5scwaZJIXZauRfolzo+Ajx7uDZnBbKlThk1s+5mkg3w6NzoM6CHGhJgA6jjr8sVfpzGUKt
NhlgpZWABdSB9ev/716XUF0e+X1DrKBHrGMqKd9XlJvd7/gVfFoDqv2Jj1FYy3FwQr2f6+9QXcA+
VKWMq7rAesBe9QQOXr/y0hrCecNXrfmnBY3Qg2Wvu08aAR34mHRbg/wRwJjy9s2kbmiIV8GpR3Wo
H24PYuQGlg7J1K7UVkOW24VDXY2B9iKBqn373m2lZcm2Q8865s2hcmHmWeqpYdjQ2EYyUrnbdFF0
yPPK/s5qFuKUuN3CkfvR6v4ZEVMCLkgXRVlucKEtZHVg8H2NWD0hoo3U3iMlkEOz2nOfg8pFHGZD
m0D6dlE86rP2fdTmb5ObDyzXwnZptVN4pWkmWeFY7uiL83I+nZkcCjI7+lkadBuaAf1KXzuO2K5W
zOwGtOjBftRO1Rt38UKNp6nC4EXixLXVVsw3AVeeIG6ci1cIZhDJ5I8uN8LY7NQqzE5ryjvURAdC
mU6ttbBsyFmTOx+qBqvN8YVa4QNXMVzaz5xHqLtkR5rKrena7ACdNnJFkZ6KKyjrpvPh5v0hz4kk
LeIqhylh4uWbF7PApTe9JcjBnGmPcJIYtp2d7dqf8fTzLfbam3hQF5qhYOYe6tCIi6eMlGLYfcme
d5YSG73e9KbrebgCgxoypuZqwKcf9+t/9sGHEQ/COHMlshhTErRmiW/4J005jBhN91R3iJLNWgKw
RvBSotRt6DAB5XU8aU74ez1sYvWT3CwNDo2uGxNDqm0fcU1bCf28N0HXNuGJoOHjw6/Pdpl9cGI5
j0ozyNjPhQEfRyO70whSchMgsTjoKM3SO/0M7H41mbcN33lvEHgitzTRMjLw2EZgcP6eRRArpKvI
j5H36lDrDtsM4DC+HY0HYAjxZVsuNzMRGuQrD7h5fOARWatjETlv37qynMvwie2R9C3BoYXYPsYs
y2RSQArj93LKM+gzQVqEfmx6u9Pk3ESRy7qt+IC7IHtCHX76NrqOtWYmZwLC6gbagih6VXLS0HTk
614uo1Z4RSv+ZnQbdeM6FV9QZummyunPhBcvDCmFcER1TYilrzLS6ts11QotFzgJAFW9hgj5C5Hl
qcWX3mCvOTfnrNMkWbDkTY6HY0r+HloNkzugVll+SANcCzVIu3HOfl4dzW05sD0de7soKnh75Akh
R8zMUL2NWosV/vE1ijS7Yskd0/xIl2S511zv7j5COseQjwGKmA9Ef75kGkUbKlWzu+zrdUdJzhqc
DqiNdKl7CbQ6AaJ2Pe0G7icoENjpDnJ4OQgc19udsPapQxEs5fetuznGHQRmwO3euoAnjdMVAXY9
ZQJGlaIZep+ofGNbySOJ9yfWbUnl5zfQdnEN0+/uI4llOBmnHG7U7oanOIbuzyP5OUxXiAXRTm9z
WiH1/sVs2ocRGbyox4iqXIj74HS6GWitdsrriFpnI9vyZcNkfSVtK9kV/mOmQdwrHNWoCQ1ITYiW
FPmq+gR7vvFCr9EkUTVXUab7AikmMksxT5UZBPwvWXosK4mxaSf9TCyOwCZDCXNqWvlmHngjTXWs
gCCtOg4cnWXWfK2L+53x0p3R9UyCaj2qPYk+rmexhqT6vJt6g1/BLbKBFn3HAHw9gdyv75MdRrKg
9Z9arjckjzaMAbCj1+6FMf99N200vmQ0Z5k5kIFnaUeAZWGuI0uHMqNJZNtqJDZQvqpDxQbXih1l
KO1MIVABVGX67V6zhmtrnsMOm1WzLdDCwKKUaROAaBNRGIExuvgWcL6d4wKOBeW9JD329d4bE8VJ
Pp10u1Xusl3B35DSFTvm2ZFWVnTpFbN+N9jE7t8utmsijQSFOEqAnyku+0MHi3Q62bF6foIxLoEo
kr/5EqggbvfNKJBqRYNV2nSDrgGRJ5nSPv8vc7rbTwhXpvXwrLs6htN48EfVl0rC1CW++gZH+4Tj
MlI/pdNZeDFRcjnOcWQihuBtFRxPc/ClxUjjtF/ddbJOUnp5k9Ikbm3CXV8GGNGwlsviOWmvvFaq
jmHohFKIBjMIqkHxJZCibNpraTCkdnSgAzHXbLfOQFAY8vjfj8i3/VycdsKlMprgDz22Ma0PVA/U
5KR9Afgp5iv5RLQTU8Li9ftkLIcFaQESP0qG9pz1r7c/ZUVPhvtQdeP7pV6N+bL9wlf1ETvd3I6d
unqt+5j9etNE6XqNiyJv6ugem3Pj6oYrBi9hp4irI3T5EssitVyTg6R94099uGyOHYr3Que+koFo
Mz3qi1+LZ0mLA0JcONg3JxyKICCyG/CiKAsYIauIG8YG6mNA2YaWXzeGEBoxQ3SxcW4X1taymiJM
iESr/d0zupbrfe/jJ9bJD73k+qOxYLt2GguqYILAJvtQCz277dvY9GWlYIBmbqVHbzeBL3gYw6wx
mkWjQzDUyEspCjeGuBmnlojI2cTV97NAT34TlB9jGkjbIIUBMWXj4cJlpoTo1tJ3Kr5BUkA9sE16
/phKNcmZg93fauf0BPZxYVh2U+7Xb/cCKijkPFPUd3T9d1/Htfu4wCVdlNiHzaDM9edF8r08Z8JE
7UONcdIznS6dCg/NcNQ+AD3ija7OjZjk5zIvK4xwz5bvNiBlgAdqXv5Ofx6dgmYEGzzRH20ZarmF
OywruRmthVkKQdHFukKMFdYRM8DQBnoMlaHoNfcJfA9+JMM0lycQ5pL0toBFS0AFjS4hMtVethIv
y3XOTcsvO71wWqBieVlknlfwVc0+pWBzdGqieox9dURoBnjrQXu6wKmVEZnRy6J5kouTA0wolouV
YMrHjw7u16MnBE2Oi8OKS4QiElJB2GctjJTSHQEOwBSvpPp0Feq6tX4zuyeqTlB502GroDOpFw9N
lMz2+YV6qW9wp0mO/ZQtTxe+FpR9vNrlUrLHnz26A51fuGjAGeRmOPBnvIjpJPS+EyN3/VSa5tIG
WH5Mj6e3avMJodO0kVZ98gX6NkbuIlqc7/+6gIW8vyxmEz7+KsFzeM7u2BbJZ11zZwns8Ai98+6Q
XYT0z6U+3qPfr4Wk+MNr4Ve2gZwuR/JdK7F324Ea9vgB/0U+v0WIhpHsIBSzvS5ty4U4RLrnWDNl
Tb+V7pB9KMVmzDdhBLbpKcfSmHGAJKmsnZ+RfgLwcZv1PpV+oiZRmJpjvXEn2OKApl65/db8wixs
EHfTN7AgY1gpeiypJU6NLWRVWfyf9R/vnnf7eR1RHDlMvf2aoqvXe9rqyMFBkTz++QNK8sXkuwIm
kcqrZUAj5b5x9QRlAcmwKlu+W3gUNngqawX/AKehlwk09pjykQB86rcz5LFEVK+BZNoxiXGIlYU2
gqmM7Z6AI/xInoFRpH7rtHRRxQyCMNzBenG1TxhBZVwkFVfresOCqecGzanNCL0PQLvG16nuAjYQ
FQ1yApxMRwwxhCjNXV2hssBZ8l++ZkRuv4X1TfV0QsEhaaXP1NW2hpYglZDoytJcZZrO9lmAtV2m
+um0f1ofeewmYaCVtx3ejtrt03Q5GBfEGRWDncj00dwGYBPz5ETQYFWobJp1CZQ7rgStdpbMRNPe
c2TXfkM/2UdbptX9p0gyl3dWnLBS4gukoe/1/xIO1Ht+hN27ZOpJ0LC4PcLqObPdzlkeh1nKW0Lr
yX7s18DQq4ElFa534WwHw7dBLQjbpFHynfdEsem9urwP/5+Z0RBb2/RQ3v0qTivruNFsmbDHJ6f3
Awe3ph/R25xt8izp1f80dL+1ZyXjXHelxGqPYgWNQSee5fjrucSqEFnW9v3aou5wJQYTv7r6QPOf
macUirKO194g4tYtO4kr9cq1xlUBM4b93a3XhXQPPynU2bQ9+dTAjFbGBPLnVggCthEDINvgVzis
rOO9gXDSkKXeQxqywuAIk2lhmyObt79+nC2DuKC82KdJryfxZWMdNKs3F7zt/YzIz6Je92hlWSZ5
gVvn1eD3rv/ot+8pNRbhMN2qsiTDnwIQPs8EqaVkNW+XpcSeYHn3pJQHD2OP+fsZEYYC09545uAP
jBeV2bYOoWIPILtZEGwW3QFANM/inlqu73v7gztKwoC0+iAEWDlGd3WvzzoKzhfJr6vyboUZegTe
U+TBxek0NktBZLHTjOtZNClq5HDLopBoeROzO5OvD+DLydEpzq5Amt5lK5MSDm0tdC/V+EG48PPD
HsmTV3EMur2YPDr1rgGzFqwfCdaP0WxAZcj3xn1coWkzbfCqmohfYfZwzoCo4fM8u1dblnXrqIpL
OEpKQs2N37K5jcxk/fkOJfZtmQL9pWW474d2Vibtnf1aQanMTrnvFVH3P4Py+1wkL8bTrdDTgKWt
5ihIF4h9OhbZMWJnpdF40G5zEvZNis3slrQo4B4s3UtdTsLbBHYJYn6a10PxHFoTI7NzWsiFtuil
BYkUZ8SCqtEyk0TEazfvHyxGr5/3ki/XHZ2OjYHIj50Ca2pgD5Uoi9+3Cb3VuSUgszW5LS59T8+q
Ks7Aw8saUjT34KZhzo1q/oMT0+tlernn2ho0htAeEDLtKISnbHS3iouCEIpQtbeLYkLdIQGZzIov
sxmXzLJVaefG1/QEuphYIaL4+YctTKqW7Iu1ylZwPYnRiPot0mm408xbp4CTZeDxRIOrYbOcr8Ce
APMWbTURMomVrTyLXRwQko/z89B0dP6yG8900umb/sJjUlwfAKt1XL14Rui2/alMilT3NbW2rb6S
tfOhWIeps32GghCrMUnsNH2jRAxKTrp2PEhanh83D1XnvXNlXMgoWhhpz1UjQ5ExlPCBympR804V
khlmAad4yNeY+J3KE426F4djNo4hFdtoCHDq4o0sLeV/qf2OF18zuzhzR1lHhMhUh3fFfjukG0vz
R88XKpv2BIT2gj9JTjmA5PCLT7/xLTkNzZRZott7mlTjM2m3o133H3H16HSk09p4x+NR3rz5FFp0
8B46I+OFwYuOpzymM7652xLNaU+J+SMHZjHMudp0dpecyfVnWzuyRNfkGcwRPumioVERvkLqO0Ox
R973MjQCShToVTO2HKcIpTqyRsUlsFUU26XCG9wV2DqjeGsiPNGF314McYg/oT2Ew9u1VKkliZvT
evhX7TPCGNWk6fW+AXFQUo5PXdYUkY670KOkhBZtLHnTBG3RD2XbevS+0OAQ6ImojtuWJsaxxbLY
d2DbKyPMKE9ICtOwK1rWOHQ7+Tv4z8xRFzQEZJNOWh6a1UDG7+oNnmGsE2GspRnA7HcKcJxioGUR
UR+KppCupoexm2ZRk1F91OuMtQh6gsB/lJV9CovgOXEBiLpCrDomAPis9dkZ+CQyEKRCzB5TTGY5
oZbf/pQtFkCWyYgQ2PaaNoKilb3dcwNRC9lqXIrME4SwCbT5DWyQMmuEgvZ7IxbHmvb0+XYyvt1H
dfMfHnZmpxbv2FWo4QgCa5Fi5VR/BAkHaudwvrJ4ENRDhrB1ODXPG6arovR1tAKWIY2d4KQctClp
a3PCXhbfvy0a+lKh53CyukocSnNwQ68ZeUq4xKKNFtYlD/IgTI82jlz1ORyqw3Pre1LvWSwsnU6S
fqbX3QGJhTIjOZW+xH29scIh+ho3ncZ86wQFGMoq0BFdFnL1lRbmcqRh98T/osfxTC0SCOUWMpnH
fdhJhhqZA/Qdo2Ck71GGpAAMsTuzEthvYUfJgEPdGiv8RZydBudEcF06DEyxTjzJyyQPwPddlzH6
fzUTaFXi5UuJyzWVRrpa06AgpdbvLhW8AcSeJaAFzpi1fmFwj4k3+dIyB4QVTRpbLfxI++WhpWo8
g2N/f4mrgNzWuLGKVp+rvMgAd7n72EfFmUhMJnXg4k/zVl33Wx4JfGroZK1v5O9RozEnBhAzmmne
RmNhq6HpTsVReAWzL/k8NsjzAHOVwwO4+KrlDU9fCyUuXHlv7kik1E7oqxz31BKIpfrpV1S8e3bz
Jkf7/Q/yiv31j/e+eFDuusUxJ27tS21UCFgS8d71EP3FvsFIC/ijubsZHx2VJlX1ZTYF8OHvzyuk
ZDdgUlSZL/5VcomVW8umlWEZaRxdKotPWkWOFIxVLJNaqqhIDCmEOawM65X7Dom91C58S6UkDhtw
oeXHmCilY4gBq8CaE+6LNr/VK0vyWYGZdiaIdx3zWrUR39DE3ov/yE+QZtWNX3Fj2ojzao6OroLZ
BqM0OvEcn8ir1kk3WLdp02LVVdZBV9YiuEAPfxWw4q7TS8ghPVNIGKRFN3nJxo1zBrtaswpyr+z6
68Yq/Y8omG/xAXq/sjbAjfMdUer4pAl/kO0P8kAz0wOUSzLsDlIwyq53MeiehmaCfdz5AMvxu7Zo
SIx6wSV5HcfzToblnsuPsmbl1ZwCG85fT7zMflzdcCWpokHfSTclIVc5dbx/n9CgzS3J8dJdFSsj
OTLTdmc0eiZNV78wHriV7QN9CBEn8M9wafTPqFhpO04QR1wDxPvNVZgh4be/4SkCIusNj85MmMTx
a60hsLHakVEF0TsXbcxJRpP8FFL3GOjn9eySoILUrRdMZtOUkZy0FS3k8qbSj7baAysCqn6oNHY2
D3RYw50RBLPza+RPqra0of7GSBNYUZ0jv1bcANFW7CEYEHuacSP4L8jrQIeOZEgtGmvyAR0BqXkn
imvnVX4FgJzAbLI6hjudoGaEGYkCxwHKi7nUEEujSVbMl0fwTaz8Y6GO1Ol3r7K5TQVfYCMdtleF
VkVnjTzysDNzcA6Lob4WvJD/RrSs7ZLRtTnyshAuJDZZirZx7JKzWerMdmeR4lOCJsIPYE2s0p80
shzhK4I872kLQpu94aDvNYlfayj72XE9nhfHrkw3sRHzeUTbWvI9S9Hjio3BWW2ABqB0PXX77dys
WaYItbElKlWDIJ/YhmadH32pOgwOA6G+c2rVjqmK/9ySGMVsHDhFafqcVE+0E0Tv7eIP4SqwP9WN
HwA0OGrCLkI+GGgWOXG/oo1XTv3hHwGMYQIvIo3b5yZOH5DHb+BWZxH8TU1t9ppXuSWkCvhTBjLW
W/GKQQXqtlUMXNuaaLif4W4Ww+OKvWRq8h1dr/Slk0bjwMtqDprlE8vI/G7abt5OB9XDO3XX2m4b
TiF/ynoCRQ630cMadkSZDvLLDhHT5crAzCAPkI4NX3XlK3V+iMg+rKe+ZeFOqKbIcSFUtKXyqaRO
2IGYXKkp4S/D1JaAZFBmnWaQjfgKjPEN4WbQ8ZJs6mXEr845mUiy03XlMDTqESi8KV3e7ruNedfQ
pSwL733xwwoqIUQkczb6ih4ZI4Q+i+Nghg+pNrttn+KzOMzZhAbUW7VcOSd/jFpe8ye4y3PgX3rb
jOWF2esAYNFBXVY2BZPG+XirZvFhUvh7it4o6gU4rfHABDMk3aiyQFlANxs578bG9sXUUj0pVW8U
vpyZ2GkFbGMJeT5isSVP7xOU1osEl/7GtN11oUZxASG4gsXjDEnSaVvJk7Kt/KyfuEUGoRSCE1w5
Z425sM+vcvk64+VJmf4yenyj0vWHH8N3I2QNJeAIu4IKcSLCZeTg/3gNszWyAyzRD9Gr2WTVqHgd
CedePnFXI6YcOBZF1nFSARXntHe5p/8i1PCmZzn4u3Y6IrGvahebdf3CyXl3VYtJ//bRkK3LLbzx
svUQYORXzT+1Z/An/BRpNI7ASpIoplIHyiG2EU6ZST9v/dHdWuoQRLOpba5SI8PvBlfBcrQGjiHu
jkkpfpk97KkcQvlvBu2yEkBDeTTsP4dGmDBiuudcXrELu28MGH+hRlV98RmXoIc9tXF6l+a28xqr
Wf/zq7ogc7McSiBi3joWoUUgIISOrfltYZ6IJbVfgQnoBPmO73AV3t2C2w+Bs1lrh6i2JUTczDZg
WgmqXzrcZ8zFVx6S+UOUHBXQWAphIia3ES2Eo8SC0zNjUVdm+P8jSUv7FiaqGoGWRwePvGPzUYYg
9xZiF+0D/5ABllFacEEX3qpI9bEAy0ECh50pB5+7lHOegOrOCf9xTQa+MtK4tps+N0xEEHLLZVhV
EYp424vLyYzqCnDQpayvqnebslpx7Zyoijf/R4It38CNVOMSC+zD6OZBV0yix8LmYH09qF+E0Uau
snXbtLf64jqe+oZylmWBmq9FQT75iwNgJ6qWLvA+GT73dqRyHw55Z+YmRosLgjZ5RXHVbzS1bvsA
COi4rtIvZdnKYgPFggWMjvcJ1Wg4xZ1hWCC/Pc6oQNrS/P9NUH65yCRHhmno2yLYj4FOUqT0dPYq
fbFHhIXCSNT4oFfwR34V8UEA531Qrpt5aPucUQz8sEiuqRBUyXsVa7KiRJ/yuafM62yrwVtJ5lZ0
EETX1ZI7pb3j+fJC2qMYY19y/xGOeVFVlTz+nO4MfGTVKTT1lDYvc6tDIGaLRL2qVLF72BwSNzsO
KwrxG9cuUq3+Jcedj/S+FdZIjz7r2fGmh73aV+PTvG1yWgrmxSpanv4GKt5h89osvzBpM6HXDmiZ
hHc04URH0HGYbMRzfyF0u3xma4B7zWZ7FlGFkX6ftqtbtbp+xgctsFUALxWwFuIKv2KBehKGNBBA
e7lqHPOnnGRQ+rnNntKNJ7UDI9Y4pGnlD6Vil2uw4UQb3klKFBl2rBy0f3TtpO7f3qHyI4jgTXrt
xZo92n7BTZ/ASP4a0FKrLbCAggIAuQszkMGlQ5bClZXzaqK26tBkYQAwkisU4kcIt/e76ABbESJ3
xK2h32st3UijIHceqoHnaSSETBqYshhyb6Ve52zQ5ND3Dbqko66n6tu0+D44BygV5xOtqRW6fJEZ
llGs5GTAyohGCBocj+atRH8ZMhG2ophtoBOQAlVna6LTKDB2fvLXj3J0K2io1D44w7X3LUNCPoTw
JtCPHfbIrdFfact1XMcUq5tpMI2TybLjR07fcJPHdWz0TeDdL1lV/K88EezuNfPw2migBbrYsu/T
jdffn84ICUXGo4I7lG9B0GB6noTLKSIjkNKSeoAvXaMC6jpdkVPp5/DXkFq3GqgbQrA6yAGrhnYP
YBH3g1VB9M1k+tIII7URkUze3Vt3+zvcCAZmSWok6vLhkQBkPGn15HS2UJWYif+eonxqp2KO0YkF
k7a05CeLvk4XEtW1rlQKCituOaW+ib0sCW4+bynluTb4fj+997ZApBNy1rvTbzdjUcRU8imld545
3xGjE0jnC2zeGNAngRL/jOC8oGRZfzGh0IUOkvkKz7ZvDAWrQkUfsnNaj0EDcrJ80jd9cg6Wpv5Q
PFdAOsLkRGyLltlWCG0l1oq79Bdplbnwna9h0UQ/c1CtY1DO1Yh8K5ok28a3Rlu6rv3asuKyeLzM
Js+Xw3utHVgjQpEJzQKVXJTbC20jkXpDRdTXge8pOqc/2BGFx2gPjYT02HW5QqNdP6YabqvOeR0A
iXjrMgObwS27bQTUw8ObnYSKnnOBCeiqV5uSQe6727btdT4Hu6gG84UcZtPWpAc0zDsoI/afwGeo
JGxUDVkHPCc9C5OA1NkLEipYfdlwIxTQicaExr+0jr6kXUR4kRaJp2olrRNGkd/bXPAm0iQsm56E
54bNf5WUQEPQogn6OL6WXnQg1Qrp4QZZoGWV6rdFtiJSHEwAUqIuk9z1/v13g+XApt8omDB1M0Wh
1i7G8oXFols5vJi/oKWBehEBK3jWHVMCYlRTXSramlAKw9X+/uxJTwtncrLe6nSZAj04LQq7cHB8
KHKu+E5ekRjpzzCgY6ffWr2clEpuxU7vYh29BRWd0DBOWJeNSbblND2A3tN4/uuguPh43snEbIjt
8RhxZ3LeW9icTkYT88yF66PkGh2CAXZ/wmPDygDkmDXklHcXZDw98jlblrsaZmLUvXU41On7Y8oc
AK1Lv3yKeYL/EvYPEJX7xW8naU0SUMHHaIW+OjrifWcmhOBPJN6WlMshVsSicWnBSptfhJhpYH6W
n+2IG9blJVt7+U6ianvv/aNp4fZSpu8iG3Kz/QCk+Qd+opKe1xrUdgrqyW+5zYAEA0Ag3iyJF0DO
PfVU9DgV3p9ut7VD+oAuUbSWAYu+5FUCwjRrEsva5MbIaXkURWNujI1qg50WsfksUn7JB9Rd5fJD
NzriyStuxyvftEYq2LVeO2YSzy+jSyOdDvYzOwE+NVnMuWanX2QA8BluWBGcLNwt43CfSwMKBEWL
6hqo6WkIdR1PFAiuwF+95P/N1xTYFsuyxZVWyXd2PpWwM9Hdu3+Y9hb0WJcBF9pbgnvBRCzR3T3Z
r4ss9VKuVXhgrk1OlrhHYnfKXQ2uZOrxCyuIJZfWrGEcmJ7PLb1xAN+bb2c3bOspBIHI5aDCXcNh
nIljrnQKqUxhAyXJUll31hsnLUh/5lm+JADyF+6ZChASYH54ut2J7+L6eMwamvtIY8LGRYed0ys6
f8aPMOVmixecfB9ki9TZh9UNrUYgOvf+3EeKt1uUUTokcgFOhrZvsD6xgQetgKrdgGzRWGpX9aE5
XIR8Vyanm3PeuAyT/Mh1wLdkO4VeL7zMDGkYLYY0+jhIz8auXg+y+JgC6HZegsA7iR7FRpo5Yx6Y
7TmE6Azn8D97n8D1CYJzbpUkgj8f7H1H9HjFjsRXYhuRduIoTRORAMMthX/GQD+CqzffIWDblo/C
SOsT8Bps1z33wdP8FHHMH5Ntnw3o7au+GzVxQFhg1DRA0o+Ui6z2Tuhx0LLI8lMkFr08D3Lit0AW
VABpeOeI2UrzljDor0JhDMmXQSdOGWSYGexEAIZCw8YkFMo/ieL/UsP+g48bDvI1RDOVcd+302j2
qow8AodJo2Z2Ocuj+kuC71j5464SrYglcArjGWk0bM+aAbtYNBufG6OVi8+JZufMPYDBDCZ0QKGE
JebNujtbFuQkLKj8KklsHqlWoeQC6WhpVPLpr9MWscv3QPgfhHzVhPzzb6R+SodbtmoQkJLA+qPW
vzHncQSKCnpA+Ocj4g4xS/1a9s59RDdTj3Zeza/QMU1D9/X1SYP06dTsPEeYLiXEXOmN2kYAJ1XD
MJO+Flv2aZpp5Q4TMg3f2y8b2XEQiqkIn94AR2z8LiMCRZ49xCgbWWICa5Sz5IM2YEiVGZ6YI23x
n4nPf4d2DOAai60dE18nl8wPbEcka0SMLVQhmnZXAhwgEywscVszQ228uJkP9eB4bO/lDEgrcTty
T2NgCMs6r8kb5Lg2hiCmvdzSTdK2MiU/AXBrZN7CbvYKELVRCRrw8yApS27Y8umo8EV8QlK1JQyO
8PNiNO7D7hwJDHB9WXrF9yE3MsrmaxST0SEu2qsD+3J1JNTPlT1aJbMAqnhznbLOZ8Cdm7r+MA8Y
I+EHPkrRPo4H4pPPVX8ttf8+BNZcKthAV7EumJnvPqx1RpBQBH/10qCFj4n5/ibCqywfkkFhMx5t
ANn4HIqn5kG/m1gY3+dJCcusoibgvhAYjjJxKZgue2JJwcYfZ3Wt5lcjn6dzcjAYVpoZ4pdvmjOn
Op/i2Q9V9q7dXCLHm6nKlmfFJ354dDKoE5awwgdQS7kPX59ksob2HY4RkW8E/WnlcQwxj50AJqWX
bOj+LBZw+4HomG8W2Pa6jvKeWKXRK1M9ERJpg7uONn1Q6Cd+nWm4PVLqwmBM5i2NoFg9pO2w3jMq
j8fNiyzKVoZGuVtl4uDREEloOt17I0xoUebVwJibhvkn+Ka+mH18ndh2F7dnVJzI8xBPBhBb4hKg
1mcjQWvVJvIBdDkYxqQtZTcwnxU2hTFRav5bTUYWqzAWwygBSg/vg8fVrV1wT5ZWx5dr/eZuK1KJ
lEYTnuTo6NyGQUYUPbKWcKzI8o2miU/PEmzHKH2Pus05zME2kebMNpz2DVsullVJpvZbdwUNLZ0B
FJ8pNc967HCvW3Q0AgZ2B/ILk9O+3iylHiPHeHX9Q7G9E5svVcXtXiaaGSa+SMBNz+uqTslEMXae
WBu0vNGGW08njTDvE2R+nsMw9m52EiIpLo/hSq1s6GXYYF/WMv+oIPJV/+OQblt4liG4puyOdnLF
YYzV+bSbixXdWYMnJ503cNqWnh5b28hLeNbNTVcMdGMnsoz8/eJldX8B1TlBfKM4QbD9b0vG3U9t
j8TgQ3i6S1QMfvUs5BWjYzvtLC7QRpZnm4LT/0A8P2Kkr0FtfaarphnmTqd0zffRl/0BtzGJaSrf
3dnqPhHl2aWSwwGWNZc/wyRA1+EWCvP0rdSwkspUyp8wRjRi0m9pEui3ko/kkCsBZY+c2vX/mYJZ
LEu2D0IGvsdkw1rpW5PaJ5PP4ztWLqKmieLI9GGwPu7uXsFoX2XyN+oImRZtTCfciZtycAK8cfIT
8S2RuBoRs7IfFtM9DF9lZtZ9lrdtXno1xtkXccTywvDz4owHwkU8RprfWT4h0ax0xNuogY/mo+Oa
r53VoXwlD5T2fYET52QyuBq969RhDnRhTwJwBNm6qh8CAyguTRGbeEHEwxIgOMOwMoZd/eYGXj72
0UviUt79WpLGbXBetDGlCx2d2dCnqDnACBIrcr6lS6s/Zz8qh5pwAzxzcnhIN5d3EVMJTc97zvjP
tcnBNJ0q18Zcx/dZqs1tRCXHE4wazXyfXoWuW8VP2ERmK/U1locAkWQOKFMTN6txHXD+c+/GYrmt
F09n8WFBoPenJ6fsfrtQ3gCW+h2b5sFTR4K/hD56RqknGr2HDei4Re2LzZBBpeMAy6KOKjGaDS3s
9mGJaKX481CGYcd0NUdh+IK0hIhLfeFM+vF+/BzRyHQiCzN2yasbZ5qxg1H9rPo7FUosE3JcCquR
EsO0R0nK4/Dv9tmZOGlSgZSlk4KdONsodM0GUk9T5HYrqE/gR/dIgLkdjf60jdkagFaeYoJVokIO
/+12orzy20yBmZhh/2RIIkBlJg2pyfS8sleV4cgHKcLb+27IEVbfJuYXG3kcaoI/rtjCkMVGFzqe
JFZeOGb6E/K8nv2V8zH0A3nBFa514oT1QbVnqT830DH13xMps96Lznxa3Sj8ww4QxNyc9CSwXLE9
yEmS4+zX9VFkuM2t0nvI+g12IzKI42rPBgQmM39PxpPSstB3N1fr1t9xNGWNE6iSS4kGB4PJ95ar
dZMzVO7k/o+wG/3Jhd1LyQVyvZVYAeC1DVldrIbmyLLKPBNdgdCztpB6ty651lPFq5UGAvPkA1yB
j18f0wFcCGhb91uD5p/m5trDBq0WzYxfTOrJFizCXsc8csONxjsU/OgY/bT14Wjp+vPGvZBX6Y6G
OUgwPu18aVwIbfnWBefKqUxHCfPC6DVAEmgxyeFY7sgjtISsWk/wa3/S53pvoSLzODNTywzA8A5D
3M96m6E9F09IK0KcNSLdmAawE6Q8aKHx8in3BAwSlfo+J8lCSzyQrmdOfWYG485jD5fTlybUCzVn
niv+aGIzSnlh//XxdPHW0Xz1f8GWdGRf5EViKchKOiX5meAsPhyASI75VPtPVMVRk8mmK8TMr+Yo
Q8yoNm2hQ83YCIsoVcsFlibU6NtjUl4Dxj0H/auO9wSrVysRGQhHzJkUPOICBthwqewhhrTHDXYS
iJtqfLWOgkX/PmsTmhhaDR/umafer7BOVjOG0wqkYG8UyTdozX6CwUXbHd/uuBY21mDzY2ZFaZfh
Ts8IIp260ikF9jdPvwXyZKC9bFSBRYDGRjk0DqlEn5qmz7FJBVpvAbL+Gyfn3/LBj6+P0/AejCeY
0jxBRgx+LzBbdApQ8idY9A6nZZc8ovz7cfgEpxzE4QXz888bKVQyUNMt+xRBtSxIw5FdD+v8Skeh
zXyP0Es1a6pgukW5Si9jpI6MLzCmThzoarSztak2Oz03GxPRgRPdBHQ831RA3wCs1pMu4U7SpDsh
t4if8bLeNRrXHK72JMrHjtWxHePgJMMgyXgLh1u1OrevDAdxIDzIympNndZINSKg7bWy52j0yoaG
RdF2z+AotXVd4awzWZL6iYLTkdOkr1GQWNuHOxUNDjR3ZTwdUbu0TmAK0Fpx5W9JmygqtsZS+kus
7gIcW4tNxYsFaQilTuiZfBXts3ZF03QSyfPfYzJb2EkGCWzawyC6HbPEIVObcHbqdOfDx1Viy9ib
hTrmDtFihdO9kP/ExtuRZFIsSwnxfHGY9CeHo7QvOUk16qt93FbfDG3LhTS+TJXVGDTSl2WUuBr6
/EX8fk0AJv1KvXOdlsO85n1rPqpisLsDeuFPJngJP7QaIz7ypMHS9IMLbKvY3FjNyjRJ8JGtzc8y
Dp+EAWptGz+fuiP0fhoYwHOxiwv+6uMeIP1JkqLM7meV86tGDW0i95O2kSLWgCN/sMoId/HXCLHj
+TdmieI0GMxHfjXfrdBTeRUWyitFPUnElT6/Q9Dayw5hyf2nhjJHSqLmVT0gNIgZdmkK5RkaImuB
RoTTaoOCWrmTrPb9lj/cSZaQBEeRYWBBVe42rtKpLlEImKxLa+zjGq/Ity/dJH/C9s8TchSr9sf2
OlKuFFNeR+0Xh/Nh+cKihFs/klXOZ6UWUHth7u/0jpKXyc+XZjkMry8It6BEpvGsH42wxrJxYFR2
iTdBqq0Bu2tItlQHXqNSEGvWY/+ue/jl4UQbeDtSH8kjFGzSybacyYglK+Ej4haMrFiIwceYBnyN
5FEhZXVW+O6xaHcznngWsBcObwE3piCW5IYrbXFIV9nrsVY7H8kMGaU0cZDfoqy6UN4+I/osixZP
Pv6H+sm5djXKSEhPZ5ykzcHHDqehHENkhaRnz2jIc/enYtwW8ApouiXFtdnsC1wBAfCcoqlJ+U2W
YTh7OoUbNNynwoDAM6PHMEGLP425Du2toWiqMyYWJgD7CTeXuU6ymyzcBmryBGx4rTf4I8uwkBrs
0+GkzId2M7DgTjNrLsOa5PBSni+CWNkdnRqiz75UhvytfTv3ekvTzdEDoQ1M0+Rdd7dztYF+O4E9
2cZzhvjyUHryOdBn574QhqwMTClGOiTlpr/x1nPkqH+PX2DYi7Yfa72YG6nhuuO6MoocWYPv4cuf
/oqJ4XmxPg7ABeiI6qDV8BlTC5hFmyz12qCGdCPC5BKZcklHb0AXY/H47wZRGMaNiXMHnqTw1MEo
qlQXjfssHmQcJkNOztetUDTR6g4YYjDrupfg88mXFhpjLYJkG8GeQcnNekKR+UOsWXJztoz1PrR+
IDeE5f0LzeCceTM7XXTorf7A2eJWBqIPe+b1wVISjSocyk3Timhgsph4spyCrSBCdGoJDS4sL9fQ
ic2EtDshkTzCUUK90pZ8bbRinqUqs9bN7IygDjG7o+GdJ3w/BQosfDgMML6pTkKl1lEuJ4STaTJT
WMWWvWWh+xHMoj/ouaAAisZgo3ZWnnYiWPL2rnTIsflYgYSvaq6f//cGuQUan3v/0gub5+b5Dxjo
479++2FIU5G8DK06eRE+0TcSAQ1SyDyODmTt5L+YxoqwhVpt0yF0MBPb3GnepjlwsYwrS4zGVYh5
9f+mxGNCGgtq+LXY/l4g2b4XqDffOOhbWgXbw6clBDdxubufVw6+dV6CAXYaKv0c7RYt8pebVQI3
LI2nF00v9hE2UzL9/6IOetWHKHFQqnhW2PkxIUzQzsDbnfIGZJWsWPJAUmT3P7ixPF6N+inmz7aL
78DQpNUrT7l+A70L2ohR5di9kyKvRMnrxxf+4mNPgIhD0dZALpCMRPSKvIfPuT7NyKqd00Nts6+k
NEn5prPTGoPVnN8PbCr7q84DBcx6Jd3lAXZ11POnNCS6kHw//h3d5aDkbb8Y2OYdksC8JJQM2mjF
cAV+i1s4HHlTgS9wB+jo6MCjEyjYEhdZ2YxjTE3fFAnO+4VMi3e+J+o9puzpge+Au4HJ4dLUUlhp
jc7CDeq5evcaBZTOVE765x06mKICfmfyCbLkSOkedzQ6aEeMUBDfv2jFlPGaBKzYJsyuIUc8IMwf
kc5JKTcfLFkLZlI6FiNybNmXU72tFKpHoYNoVchgLYNT30z3s9365k/DphZTSOXAExy2Si9hrBmj
jDa7cK4vyTebDf8Be9WMy6m8iP7vj9ANRRpfSbRkdAgup53sCJMOsWDx8JZJSQOdAvQlaTP81ORz
YZTm059kf+8zeS8j8Kj8VCzelwzv61X6qtLItOET13p6MTOCx3KzhHrPZzoKafJUQiTyoArSWplN
jCRmw2N9nzmI3hHxjWnGPqQQwwzO9HZ/pA1e8JKpoFWAmeTiClKqJNoUY7Fw4be6prlbKQ3h0gHt
IxmJla1zQq+2BviB9RO37CxWzvJqjVZCNwO3Rpos4FXiMXAtPVgEXjpteXJObqNBbhNlygFngC6R
1udROmUkMVnHEv3zjyqFLQpnX4rd6GaB4yFJjDXKAIClNbuPNQXhxTZXt1Vx7/3WkZRvgzGkWMWw
IFNI6yDFqs7ByqvN7oY6g+QXEpv2OftpyRhSb4ts7s0Nm+MLlGwUCer9gTqCVtpozIZIyKf5FEHR
xVPFyQdWA/UWPOFZwFLZrZmJUx4K1WXwXg9/IKwFt/QrD47jOnDJ7DhxLxA7ts9l2EFyzeEMLOk6
AkF15AWxPyin6O87UpzHwgPuoQ6J6oVgW3UHDVhfrR4jkFlEYlGCeCRVV3mgtGWMvgwFKFFbK0Ud
pkbzJmyd9WRnht/XwJiLxURWT7lAinEXWywvYudUaT8zG0WX2FsL8Owp0t+2ali4b9TEmBb+E/Ne
Za8PS7nVq/o/IZvsAYwEXF5l6IG39LeBvgDKUmvCn87rxG2xWd+D6evVcdD3my6I1BpdzvtIR7MD
DS9trfZjIHGgCr2Ihj8FZoqBvF2staKCvWRLguf2Dl9USToJdn2484WYVFVvNQMzYmJL0jjQC9+8
9WCUihzPBUApaaIdjkzdNSCvVXdu+LmQWIJEjoiF+wSWBzlIDy5xSHnMkddxhrluNmcMyPA2tQZK
HVw/P7pCDAB8C+l8FeghmknCj2eu+wetySZ3ViZCnL3+vu70ZfBn5bov8PJxUVhJ5jSFNuFL2c93
OFBW7EmbwTP44TDgr7ycZt7NFvXmD0QO7ZCEvvKJZS2CQXvMRZ/JQ9pFP6yoK5EVWi97hDZM1IFx
OIHGMKP2S2CCUJLMPOPxWzNBh8cKx4iPmhhwEecNsXR6jEh85tQtUQZPfvvhjDfcwSgSaUrD3Pl8
qwhpL83wNBP7GHZrG0fGlONBXZ8BHGFp2reO5fHtlI6oxD1TK297AwXLqceGO1XFtYvmI3xu1QE1
Xw4N4Nx7u7Je/2VvUz2fGhLegX2rlEysoehx11SytNxaYk37nIxdAqFp/pgI3oaT0CDrbWmusTAC
O+8lZ23ueGyEpIE3EOH66QRmSPkG3KXSdNnj33fuJ8k+w+9I7TlQjiOXW9cp2w7Pw4ixox7ZJ4Np
Bw5OYNn9nSXfL7AMhGUvaQ7m0UJO/dcPu4Y6CVf86XhPCYlTTcEytK70yOhM93YZ4TE91xMVgrSb
QFyxZpjHy+LfoxcEdi7vOhmZgoBajd011pAcATrFof5Q5OfdolTrKBU3XWekw/20N11kpIrsPDD6
R5awfzwUURcRFVCVmpvMXt0PxbKZwCd5cAzihE95CrRmjxHhsLeaiFdaOopUDftuzuhxAsE7+Jsm
jQcYTlWQrx9aiTWWG1ktmwnNODPfS0vpskFPfoqjvhANheFYLppI2yB17vcoLEUJ6gK947SI/Zfz
ogQ75t++cG4v48UpROSSBpjDFhZhXVn+/wirbfi+Jx5hPH1HvmVRWyJBNvYwRdWuTeW/5oBfl+CM
1OEmpYooMcXpeJcSO4+7UiExt/1ZmVhCF/5FdhvLSQeYevwqUUfuu4HfGTJ63uVCU+5okd37a8BP
qMH13CgomtgLzsv7Ia1nNHK4i/6TgVX8W0JRQapK8G8PQyv+I3CqdGJPDzogoq2T342BqY9i5wMI
eqGR1rvwqK3aP9abaAf89t9ejEkpe2h3WJqziVrLGxi+5l3060IZ6SmW/M/WiFAhSpBvnq0POYIQ
V+0CiVlmadhWZIQD8fSPbizkfN6zv9UTivGVkiZVbWvkmvA3XXRVU7G764PwfP0Nnsr92W6XWZN6
1JAHXSdzRMvyFpITM6d4Qz1CHfJjC5+AWMwTa0KW67pyg+NzhVkCmD510YCMzRPZFQ6jMNF7UBoH
DkbwKp4h2lLaf7fhSNtGTHO+Zznt8u2yjj+cthOXfTgOmUz9GtvVesnw5hHNQ+hWdxmtPjpNHYsm
nNnHKLN/IdlH/SqSu4akDFbFnXvWy8I2ywLCfKdCgVyzuNa2Su3pN2wglHgJoh6WqABP3OhvKFY/
b5YE7StzK8fWaq2s7GLB3Ago7ZTk27r/cVbuG3AHcTI+gAQOo1I/qRomi1a2pTEFu2HcpSFQUUyr
Whk5uu0VwmCQf2TtgoPUg0RqVvifQqnO2wBoc9V6DGjcL2CKaElHJ/LqWYA48h3c1WUi1Cbo8jSU
U5optj1FrcKZe1fRJiHOKgSS+1rZtJr8WFvZb87XSqwrW2OvWVm5qmQKiNh6ymDAfzUf+CCIyH/d
oKmZ9aE0ZP6ioBQ2rW2jTrqDKqB/3KO18cHxfQbchX5lUEI6R/pNEdr4RuflTd1MOPvuHfbupmX/
+HFdHKblyPldNqrK8NsfSRNilgyyylM0uWUE5lCP2PAvzLL5zwAVOb7OAWIM4C2MQVR7U64viKLs
14PlafF9knl78zy8tQY+GnNAvbpzZlJb9YL7M2iSQcHTqE8h+IZsz51ZgU3gMFOs2KYw7TJA29HX
mg43dPz/zaJPvwRQYNl5ply7mo3hpTUw+DsuLrtzk5GQujXsMO3T/2YOJ2Z5kWrU8/gqrQxFqFcK
f3sVZnXdYCt6raRuyp8J1PzDQIrHsvzxe80NWsfMgQS6JUA+OieErHTtQibW/9yX0FBZ5BV+JvwZ
+tWzWIH7RfPmFeKNaqmrbhsRyn3/ubO1+yUhmqb4l1MUmtogX5cTpthbpsQkhyI+he0uuq3ztpjp
72rSFfrVPqf24mEIzI+luJmemoP47VRlAlp3wgGPD2G/yjTyrwwGuZWR6CCoSIWcgiLa2LRLnECH
LbRaAeyxwWxEmPjepkUzKn3OFIin58pkHl3KxenJcjgBLQMtQUICiElLvghza9HHQnhLxZCFpR16
Lk3bg4P4aZNh6yuC4EaF0cAbDC28M6yJY6ZnhmYUEd6jKO0yJk0N8AXbo2240V4Lk5FKMwyAf/DQ
WyH8ItzTqKRQEriPlH10XhRTKwK8KYOty9v3LcHjMpKyjcmwInLnBdfzGg1n/tJbbws/5+KLdhp7
Wvc85Pzx5zx33L/Ovt2M1i853IhX50upjlamD04k0RiDw9C2hHp9qx6whQ1BSX0PwleRmX79gl6d
2n3W7uzBvMPDBvcQpoKvMnuwMoJYJOh2W2Hr5b9y2sTfOZ76yCpMTX3Fa+Mv91ichysr9hEh8had
B5eiVdvQl0iccnUohB7nQ3gfkp2FbmFTd1Dvugvrfr2AE4wgxPRtc0pvU1ReMy+M1vkLahlq2qug
UWic+4oJJqCzoCZQ5MakcHRuAJOIuVKtMP1LsAKoYlEL1Y7n2sSZJA3HlHGFTrmC9eRdSFp56rGp
o32zexv7PaZxriFo39R+Cgh1+bcLrixdP8EZFnP1T81rJAMuyVcKnbWL966id4wpGmBRwLibqv+6
/R+LH6ujmz6TZj34oMc1wF6jeelsb57H8poVRAs8hvS9WqZnwmHaP4RmmTBK4Bog7go9SU6KmMjW
pdMR6M7kLcOxcn38W4tFVbdc7jRYsYEtGz2oEjfi+i3Wv8AaMOVRudDGSs1Qdig8hCE0th2hsE3w
iYSbIrbruVaQxr5n3jqJDDhXinikPYyl401h54so9CCaZw79s/w/vCuILRlKdbOGZYMaoDnmjZlO
sOl7oo6Qkh+hAqk954rysmzD8eRblo1azNHRyKzReqGyVEYi08yiNTa30sdp0XhHmZmGOKAmkN85
EscMNLJcJTsArJTvBCE4g8ExPSxydAiKl24ONEvzvLLDCjksSO0vSYR9powGTXemKi9yUnMD7/sA
ypXDwJW6blDG+Hk7UCQ5o7It4MkqZOzEb2RFc/klG4JrV2YDNkmk2NLdFktC3+EyO7nw4GO9tcl0
JNzj0RfvKdw7VW1WKpSriYSEqNpCyjkBnmUpzp0rn70HuZ6UJlf9C4Y5dVOFGl0AU57lKQKxCJI/
Hc4YMMmGWpuWvM4giC1l2ixZAJVWYzfp5VVpBv1L/WLrBOe1l3ZAq4FOZd+1PcjOOi1mKyIoaEHW
Twlo7lNRIAJoWyf8OI/toPC7eihz+uABq8yUpIMSsasI6W1j+5CioMSmuMx88/oAozCkw7Yteg1z
jdk29zDx1ZUPQTwfhVbUDkKRTR98q81RhlzddAdn2SYkEEMa2Y0Y1ugTQG8RNLcwl6rm9uj0a9/8
BdkOTw3REi9+OVRhdIRvbgrMqjbdUb3P58bF7MjQe9/kOHgMk61RaAAUmWXeMvTODjyk42xqzVg2
xG70BSks4aMdZBsS91VaYTkzvRa3/fDgf0B4O9xiNTX94IwikLXZltRvgVTRRi2/Gn+bBhovR/Qv
V5Aq0pZh6tJooFjqsS5qzIsn7t2bcrrxmIEiVhFRlclnGMDmNy9E49oVviD4JD4zRGatnVfhHYK7
G1P4NF4cbohblxtsdC9F+BsOGYBlgFRDY927llM6llOFHIdEorUOTiMPAJmSJEUA2AOmyQyLB8zb
Cqpz6rx8nkWNZqgA4cFFG8tvu64T0CNH3WP1L1M/k1oUcbDsSYHshhOcqiUsHB4+DuauiZuv5ktn
cOCkIl5LozNPY7ZmFLWbY1cp66z3DeHKgsT7goijJG6xrA74PxWNWYZmlyAIWkR2BucfZGBFaazn
b5NJC572Lg6G0GHWlq6PC8mVtflvKjAGQSkvwYobI68rPIcpIIS3N598XN7JRPUaBm/xgZ9wuzP2
O3vfzTYpOjqEIZOqh8GU5IWiWSek+DrEw2jd9XoKg1wIkdmcxx4TU0H29Yo0zkq5Pg/+J9RRuwUh
FgKuA0nWQUqllaBQFCbYcQbroJtEUhx2aZS/AtZY6YZSRoGwxpCp1k7dcQR0z+A1zt1jOpcJ7Tdv
TNH617bKOyFvCqeXdtqtCVi3uiSfWhUYj+1sKXuSbalxF0yOHjHw4bFXMroaEBOSel7aHYTR+bnO
Joql8FIg1nOHlSmGzr57uruyxb4p/z+uMZhUakZZS7U/shY8jV+lbN93y8bhO7ent6tRWdKdJRNy
d+ez+HMfe3P6gcMxou2h3mPT4tsFW2OPz0zSBm8eFoEVyd5UpA58C+zesH0xOHsBTT358zeolie/
CgsDGJF9JjGv56Tk903rIDRFTGDRonGNQq+1ET37CZofCfxUDUKwzxq9CAkiES2BnYeG+D6MqLKU
rKnlXPmfxTDcZJuMj5Gn38XUwf3JTt6RIgV8CEqMnnnJ1kU/cigB6aS+wwRO1bCPjVNWBJLgSjkh
mwsTKqjq0P1XQRcbNQryfnWXx2kTvIes9wAwkmf5/TxEZV4LtjiO63hn8C7esEgdHdsyryfKhbEu
Cm6bjFel2anMS8GO6/n1omclcoRaBclrvVFL9dWRuAFydRDGu8f8rKp9hmfrAaE9I1NysXIPKREt
V7yi60o+OG6iWzlDPRG7h+0HaIMrMDmX0ECwRQ/rHl0OxacleUEmgfpiZz4ofX4stwcjinjk9T7J
kAmbJktXEjoQ2GtEmQnjDTdtkstjYQL48c9fP3cbh39R0HHHzCIWxl5smdi+nfdrZYuZqZEj6dKg
IftOf2TLO/Rt0qr4TJV+mASabQX+PJNRDkKL7UNMbwt5bfFfnjIQxn6FqSXoLq0tAyGMFWIDiTID
TNxr1vy131S9imcnYVcbTyqaeodsxRQYn369l5/Juxy+//Ief5aBRmWBNh5avidCVA6xbmezkoLl
YzV2JcUTX/nM9g5hVAfunGbc20u+PkWAPgwwAP2bicLImpc+GgmpiWPw3JB5W+88JOc6RMdwH5Cu
zYVJNwpzsyc/kkvjefUuRLQICTZg4mUj5IDSctBVtXR5TXhoZhE50Wt4Hss3vEAo9r7Z0yd5cSGP
m4mPRjB7iVrRC6Ed6wKGSFLEzU/JcpyLXI/WJLxkhK+PFNsIVhcC8rRZMi8yQ7LCoq5igK15pp4W
qDELzbTPQsRFrY6Gsi8oHwzB4pbQAV8N546k03+MsaJewtc4xSax9hNT6AXGbSqoOWYsao4kCkbu
0+JeEXBW7BibbCPSFyj5yj0YyJNKbCZ3iTwjG8Ny+/QPne+VJ/vfSbDCcqUxwc8BfJ9jJKG4CyVt
4uV6ZIQud3j8pbIRE2riqO2YDaemlVM3N9Cx0Gz62OdK1hTnbwTqFgfM3MMA/aQ/jXMbcYfDhquZ
BMmi/4gW+T1u9ODitw3T3LjUR+RFt+UwIyU6aqjJqMd9FmoAxdQdGpuYqmOFIyMezkUywfQVGxgO
Kfxb+ZRpj4b1OH01LjVYMkCR05XTDB+dzKzkhqdf5tkmhhfW7v83HTRn8cNeRsfHNhE/su0wLfQ3
AzHwPCozdeAoEsgSSJl5cZP3wjQYe9CV+XlkIcfFS9iqqMXqH5inxK7Q9b/snskzCY+9RX8EsVzM
zf8i1CB0IknhYoRHWqpe79gmYoADi1lC+1VVimldR3tt/znPB6sjCX1rocbEbJvn/RWwQ6mxDyVh
4p6bqA0nECtRBcjdGErdELqqUD8S9Fn0ZQ3Ii1S1KEV/umDKQuAtcXSAaRnR/lyNdn89HCWEqhej
8vv99RqKTBhRZzM9CDEmf1zPjX+nxZm5rMPCYf8TrSQf+A9smjcNO3pPWCWqoyziYSL56M6L28eL
80LPuk4GeUlzUuEWn1BiIJ51iCTT8PotGu7cAFIYiIqduVpwi5WBgvj7BLN6CZfKJmq6TFv40AzN
w+5wO3DSLhH45DdbUwYn+gOqC6Ndh6M7PT83O2qU3j74XcLSCgOqIjX3I61OFEyqkC7B3ylCKD9G
CJjyMrTGssgD9z+/KDgYJykOxBfwQIgLAdYMrvZdMfCEPWtya5+joQFQgnZrrfk1ijfYPblpdCLU
p2PB+bbJGCKN9L6QUFmsPS5XmIOhp0J+gf0KPp9Zb7We7AHTSoxFiayHzui9o1O1XTdQgoG+ps2q
DxGWmU8ESaiTz8UnJUh6ld/Ep0uV234LpBHUyhNGx+dr+ZX+427YZki53J9x5sTYpNrTFpLEWmeO
v+oD5dT2iVaHQIc8gmV/MuN7PbDdQPxDBoZe9YZf5U0V3DcjkmxV6pRegA4LXDQvMY+u6FDo4f8r
qJ/G/EKmy1XYG04E8PeoJs3K8HPHjO9Fw+FIfOOdPwWcUgi/oSMF5GJ4HmB2Dt/0qHwwDZBlHIxF
kRxqq8+3lMoKZ7jY2RxCKmSOy4wuc/r8xz/epuVKw3BafcfQXgddm/ghgYBTRsCDqWW3Jp68iFdD
lzxs8ErFyr8yCeIklyyWAPWVQGPmrtjio0J4IvOusGrkSnfIS9dmov5dvKrhvgFb5EiCCw+3CuT9
3j6Eq2VyZ9TP964cNMfVPAMRXkG/Lh1OGbX0xjiKiJ0rDZp+PhceFM1LKivRraVVuFy2FjgSDr3q
F53x8Yos3H76EIhF383FZUPjRk7PcpFQ1Cn/2BiYvvLCTwlx6wY4wT0byY+2gUmQEK4MS/klCYZY
XBKZ+iSguW9AW90At+462ifg1rftgbH4x7sFaGsAJJUp9R6324unWXGPzTAeXUvvAdJ6Ip6p1X4X
HErRwWnZsf/UZ1Swbf+oDJDtwB2UJUGsOL0ugnmXw+rBAwiXJnpcGaAZQz9OnfoQMfeOaURk1XgS
dNFhvxelPQESH+6qU8pwPS00flKAtQoG8B5bBG0W6NF/zFgH+gxk8euQr8yyOOsqkgcPTsD0QJoK
u8NDaqQacYbBuo9fs4EK2vggixYhG6TPBB5lNq1fdxqeE+a07pjSlID5ABek+AogrTkHUBVG/tjR
DtAwo32sxsp8YHsXV2GjFhhYMwHdVXHfYSp6SKsR9iNg+f1tkJQpsNqNNUlPeYOCBtQMdF3OQ0mo
STgWgPs607HNYPhdhIeKvoCtQ1jmM5Hp27DKC+pq0wIpyCxeDfBeLs575FzANPftY5pIoRcjnXeF
eOogOvkVqCE1ZY1SYP18LF6wpZLozOS4LAAGqyGCoCiAL9L3odYLC3qZMch+peJiZ6WacxsAX7ml
UmkUEiPXiaxxfQRrFjLmxCPf1QYF9a6cdLLeumrseAkCtEECQNs5krClV7cwJudWn0Zo1CMo/9f2
o6kS5gOaUCjpywg7FiWbI5cfbeM8FUt3jouvVT1vJYdW0raKOOndNEgo0d4YG7ufIVuGWqY/+nYU
k6HepwO23oY5a7Acy83rdM9AVk/3IKp8gn53CPOQCqrspT4wObSQaf2MYng+Ti5QptSqi3Bkg/L6
28JxMpFf/H7v++A0M3Fogj5WKiTpLrFmjp7PGDb+F0qKMcri2c/lhgabdksN22sykl+acCZ7yrXh
EmgyqSJTLgFhs9binQvUhhISjOFsmGGhQUYnSfWVSz6JvcZHgphkHnPBfDSG9haVZL4FKVPQMbo8
bECwApCNZ9p4tpjeMejf+yiUWnsudpO19Irf4/cGs3pmFjKRzpaInT9kFmERcOkgWKjkYEi+fqbe
T4A4EQBn2lM2XkpNe5j0tp00DAU2iuUgyR+RyV4iMV0chIcc11xjeGojpufJyTdEATlJGK6SxIkd
yICj00rkZZWzkyfsQC4o8YhMstxTPCpoea+KUHAIAacFFisJYIHUDfepV9YabUs8wt2v1sdRwAW2
YqXhW2HWdUmKGqhdifgo1vfxH3+vpdiHVdhgAougfwRMC5vOvETBeqz5CYt2mK0rofyIbCc+wjI1
i85uhBKEqF/8/dJTxS/c0ZMFnaoV4bKUMA/Y0Wfp8RzvvySp76q64+SV3StfspusjE4lJCLNNO8I
/zOqol4Pex13owg++4VKlVknkQyvUk11K5ZlDe47wD5CWuQyUxAeHF9BWmGqJISVOXMZra9E0hxs
moX8ehoF1aWepJIBVCqoojxyroHTpR1HDft4LGWeGopWh4pwQV/+179Aw3bXGk89ibjlpUPpafeG
jpRsEqNGpkbm+589lFU8QPRD3RLCDfHKXZhkxC28i4crN5LJ1sBILr94ZFWy2n4sRDr+xATORLe9
4MfguLOcEyp1bOsniDA9X+4EQE8uT9LvXVZ1Y7dyS4qCF7mYByqjOK52gEi07sPZak6XBdqOxNU7
rw/RRHDM6gAHSEduFd+yPvboCLvzckuD1OETzF3nZ45oBpa0kOILmo9e0aNnrLNLUkLzopEIhsAY
UyuTWVJabj9bGQPmEdWjAiAQNZ4eymjWsXDVTFuOjkC9Vw7y2vdglF5ALNqVRtOpoVaGAfkE30Nz
PCQrzuwHgWeLwUcNxyRV35NcK2L4+p2swWr7PgMRnOSj139Ca/dx3tyaPR0uGe0avykOYl2iOy3B
w8i3pryd4C9WR0WRTpVrVTt5fOTv42hOgC+pouo7C6ISaITrPhY0JKt12UjjYg3T51nTLmouyu5d
Dnmgn3zEjnj9JDLGO7VvEXpR5yJUz8Imz9aZpwxHGYmz4OXBabiugtTyJR7BINlw/bJ/NiZtFWG6
3pH0RnvYQXe7nNZSDQkSm2x/ZEzNb+Epm31lpV8i2f+R1VaQ/cOubvBS5LCqenld0C8AnFCDsVdK
HiN5lGdHAOKb7HMq1BvJwhCQ+6lsnM/DPty+UyA1sjUZ5wzfnbtB8IUbw2Qf8G+zVQAwRELGOAjx
l8cP8d7spCtUUrkz2S/r0gP/8Lxoe8ijsL0G69x+xDuUdbhmf4VGykcm3eJKUL7ken/QZODTpKgY
PwBN5iH94Shmse+pdJSqVSnhzYkjG1rhtTi3eZa+g5T9vfzCsNf0TVa1hLw+DKjifLZlGRGYTFqS
3/B7NkbwmQqyyvnlFRzDb3QsHQqvGGm++/cUNbxSosdRNJ/1MkzWSi3eJpYaaPiYA/m+pWnJ0YxC
/UZDtkGUdDnxcU1SFQm5d1oB9zyuQohem75FJk14Mo5AyO7T19nFqbyR9v82ScJRPhu7eDiepkQF
uHgiqwa2KWfTiV+0pXFBVWAe0T9CC0imVd94wikpS6nqEzI64+f3Zsv0rmhQu/cvQJHDUbGIjDzF
VvkPkQIu8+fbLYatKGZ7COdrK5hH18tVUxXPB+XjL1va4hF6vMesAAZm/S9XJqHi+eGFXjSXWAwf
Y2dlOW3jGslwObnRdF6nrHn+RSWgd5Zd3PuLYN51uZFeVnQMsNCTIz3OWQJonJlEu8b91fERA/qy
82uzmGxpNhLXMj47QkO/vNyrMNBUOQeCg6KsgVKvFyYRhHBDSA+ufpqJkivRUD0D3ndhzytHVC8A
TkC99Fd6lf4zG7fr0sl6iSPHmXkuq2xxC2RGoP+hHWMm+XFRONsTamWzjIJNMaMb5TRKSlJhK/mS
RZ6/jyJnpSzf8sKyRzRVEHNhtyn5vrQG6LlD1MSRJqpsMTKeopojsccG5SHQqi3JMViq62tmQYIt
MW+nHQZ7yBR20R6ba0dq8SYKxcBcrbURT3s9tFIlR5em3GIYeBU7z5wtku8RY2ifFeRFBmzQ9t4T
zsaI7QbkuNxEoN0h+iuQd/xiDSrfT1JUsv1jCTRDJQUkPJIedaSuQVbraqmSJMqxZBW/qX6exK4X
zfSS9GiS1OVMFGJ12JF7fqH91O1skgoe2YGQAPWkxcSchPyPXrQ5K8NcBYdoQINLURlhrnqlaBBQ
K5MuTedV3brpyoHASe/aFZnGHCdzZ2LwM9d4ycqRZ/oaVfag1T6AjZylJQqviWS0vqzQiPsZ/loU
p9zi3tOyvShBFx6P43Lh/wnhQ5KebKpGrPyfTKURBILEZuHOxoSfS1ephtb+RTMGBiz2yGK41RyK
fEMzyuVGX3pdbSsSPcU3MgdDxOS2nWmDbuONCmvp4BbymRckxrUsqGqH1qg7nRAsrGnp6qDVieyc
x1ptVjzo9GCpwZ5Xp+9mBh5rbQHHL4CXXzO/MGOPXq8wch2jtaQ4PIz2GzZwMdRsVzAi1w34XJzs
YExaGCfqPGD/OXTejgX0bpAj7S9jPXkOSZ+wmwrOSaajKuBZXJSHZbdJ7vedyibPc/97H0ZpOOAq
wLyv15qiut4ZI55I4zHrDkYf4f5IbEuidtnYv5MMfUaA5r9LcoUWUv9Kcdrt+Q3t5RdpoJVTwFaq
fAXmmeTzWXBkiPg5xvOQThYOTtMKXdff7Ah2fIMXdR+6BmgsGse8WM90bjSMRqQ/50THzRujM2f3
b3VngQO9Zg78XLnAwAdXSEf+UPPiwu22HCe9DzFD5T+ZG5rEx2tK6ssE1yof2v10YEJqnMTZSx56
29htoKxcy/tq/lQGcLwKzHsVpJBUs8t4o8nVerBu1+Zs9/B1y4t6fnkKHhr9tohyuZCw9kCle62s
+ZIxFL1OgO5j6BhTAEKDTTMtNYsoUWsGAA32kqGP
`protect end_protected
