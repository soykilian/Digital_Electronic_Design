`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NmVWAqENwqmr++b+2vDwDO/5hIJACqRwrf0XQZ3BiAanNgFK6Udy8IJsYu/5ZaB18xZU1dIS95oD
TEw8Us9lVQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
keay9vIlMTMToTnPzXwBOLzMo6/T7cfuq/2+qFMTtZ4+18KPY1Obp9/Wl7SIUE0SWX5KudNn19GO
ymEY85VDJAT20hYp7USdIuEUvmMmk+LdSDg2ebj3DQJ2U+h5SIMEpPByZGLr84DzpYCYmORYz7if
0bfC4O4iVpXJ0s6XvL0=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JFef4GMguYl/4wXovG0UKnYdJGiVvz1xUpme231NOhaqXrU1jO6kbs43l+Yx5Cr8lzER6+ocWyMR
N4jJV3yUzjjWF9dAyG6/9pGf/8/ajGuBcPGvkZBxp/pA+YDA506DeFQ8CAGDm6c78JXlFFpqZtNQ
VYQx07UfPDRKho8z+y0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DayeqZwDgXNQ8cHwjg9nSurKyh1M4XEh5Xp0+4YPzzXisB9PodE4Om5ut5GJn6/pxM4U3OVnuc4C
GaZfmOk50oER58mk8jIPff+oMODb9HLYz0JKMXgeKBR2ICNPQytRVM3NASvQNCFRTA0TM/RJIlUi
OA6iGZqKCOD78J23kkVrdDrwjE289WhAI3IFpThvB4Cc+1vXE1jVafj8Bpa+0YY/YmQlOBiyK2fS
pxJT2MO+NCMcRI2nlWz/Nz2sm2xgufozrvyFimLkl/SW9y0i/h/Jxva2t0CCHbepkcqPz5WcAv4V
bmUQzS4Y+NalQzbrNpB40sTUPyeV98FVPOCsBQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kYkRbeXN9gAcs5zRlte8NzSTQ5L5nUNQnO6Y/amVeB6h7JF41HZdRylNTC1lHi9GdcUxJ4V9L0PS
jeH0YFmqNjovEGgG50DagE+YNX1FKKmPVYhS9KIBpyKzAJD6T7zR9tK8gSpwTgOGEqhlLrIxDRvb
uIbkhF3frb8kJTjs3EvGyj5/g6KoCWKhpS2tM2crbW4KAU4Cqx22HHR/ZpgBh5e9H0hqkss0h3HU
lc6Mqs5pyTv2IcjWALKfeDVIpot0RnYf+52tlqGlFhxJ9zehW72fJn7vD8vZXaqZgUBbaPrJKfl1
S+jKKh7e7VdWWqKd3xvpeb0wTrWIlvcNil7SXw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RPdrjHed9ztwUJfL6qfSuAnDbsyy/LPOx0VTfms3GRxCyDktYs63DqH2bfp2HfxGoB7EKwzsOCSA
WD4U44uVA8QquXq2To0Oh2x3JBSGx6swqd6zGj7/Efyf/vHRqNCu68upjpJT0/+4KSedQT1X156t
oC9C12geXfrxXIIgZ/dTs2OCWItGOYuCAOvs3+4HxfwiNd3dwqa2OxpqY9nejLDO6+WKYrQnW5aQ
DlhaVRepa1ha839Vstpfs9zYpDWvwvYvhyoMqeGidtFs67/w4H26q0Ev3B2tqoHW2J4MRriNG6Nn
Ixc5YsGfTh857dmRE8hmt9Ghmqfy8c1KFY38MQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99632)
`protect data_block
U/wAY/cp3bb0/8tCf2l/TMaenUVg+wGlkuvAzZ5Y6XBwiFsTBacgmGRu3b2acewC6P29Am0csMmm
PPHC/23R49dfDUcqCL+8HmdXOmtJXZUk9HVGjDG4phz5F1bCSawpYfeflQSFv/TWPOB3qa3YbLiK
4ybR6YlLP5KkEd1DTt2Vr2yyu5okwJi9sDWEZ3TPDEjp8n3XJx9sYNRwWN26YRCC3owrMTtp97nZ
JTZrueIlDq8SI91Hg7MwcuEymS3UQ2pZDRxsQ+nO1hMa75P0v/pJWemL+ATqu45lyktcNllyB+ev
KjIhhRQs/lSmI2jCussG1m0Zr8merhhIn+747gsoji6DH5ounDXUZ82Z1DoC1IkzxSpYlX2qKK3Z
X+odT61UNjy8y+Z1uYk1q7wWgLDX3gm38xET1NswDBA/kYXiyxoWtPqLeBbxnTu8Xlk/k3zhdFAo
rGsyw4WxvxkJy9wNTEKwRBPF6fE6AdBuMctlCF0TLqxdcgpt0DYCPbu0M1sPzUnK3eSmySpAUPZt
7C9/ah1uzIPMqTw5MBwKwJT6FuYRu+eOyj0oox1HG4rjxHXmJlEzDp0t+FOGqZ6OeCb08tatf7EQ
gBxm9J4bXe+lx0mygiyMTHvSQ8smv9g7cN+WEAP/GoQNLcyLx7yR3HzoROBDhs1OAATUwSUGUwRD
tnhg41e9D4BpMblA/5fZrjrGvfc6rd6452m5xf0FuWyiOtpY86UdlwZfCzzkIvWVgZ9TwNcsoRnO
I+zExhB7+Sc2a5DXnX+AZXS6r4A/67/eHcZf0jib6GPoBOLkJGoLBsKGmbV77EPdVZCHuVaO02Zg
lPXcxZgRIC7CvVb61iLca8o85AvquPxsXvSKXTq4OHvjq4rUl1q/i+PIZdFnEBk5+X8fw2I6Rf5i
XyJ5XD6u3M50ZXOiZRBoIH4yaKvMRUjy6pufAo0o01O4z5vSa9jITBcyqK2ZNXo2HIo0DA4Y02nN
15VmIex/SVQGaGhnbd/lLKdV2+RhVCDsb3TLfA/7ZliE5KqWqyJh4BZ52j1nyEqLQ9zEZorgGcHl
r2r5PZnzZV0nEKqo5KHZshtnKGdKky80YLLP9Y1GyR7IVlBYQ8SHQYSKBe9qI2XpUSKkvjBfQA2S
3JZCfCuUdND4wL39KzHczDtCEpjYNgxAGGX0y3fvUjScv5ogXaAwymlSnmbl8OqaNxQUBQPkRr4V
bIeImr7BC6wEjDqQw5B3rW7tVmil4nt58K3CPhBp2SuZX+thvM2P+tAQhwkCMaCmGYbiqT5TGK3k
WFXArqzlbvBzWUf90KgrhYb8lMl7hpAExik3tGPfQALejfT+qBLM/3Z6x/XPS4sJsBXg/vTzS4Jr
Kg3gUcdbNbmvCl6dye8VO+DmUy1wft8VEM0HemnbGL0kaHK3t8zv5C/SwrWi1Mc2QFYZdQ7hc58M
7w7da/32QM3UVRDX3pjf62rxl3YpVU/mW1h1OLucUp1jvWxi1zJaLBIpTjTl5qHm7Gv0aZdDFni7
w4yDVdr7fzoj10LkWaU3qGCnTfrkzJIYCD7R8I+hVEHHcqQipgEPbdYsZQGDe3oSy8ZDacH3CCwH
7aRCpzWnoKUVIWzPRv1+AqxBU/U5h4zcFHU5rvmf5VLNIXlVhTHQHDYk3P/jkyTO31bA0EIkdKVw
x6CItesNT/DkHfuyYltZ/oKxNoUFZivcxU+8ZoMsotXyJ+xdcg9bkb4qN9W2yZBH1K8ZGuckuQS6
L/V8Q8v7lZHSeFchgZ7C1Ed6xSR0gktgIX7mRU3/Bd1WKnwFrZ1oCzw7okdQvwEjsDjkC1wliJlB
GWQ+qmYAkTArTt8OVQgnMaLcmozswKNIvgk2Dnh0Lk0HtIFNPR7g7E16hU7ZqvJ2642pVXOeCxH2
RSBb27sfV5KbKdAHtA9GxtaMF48f5ZoBaClxuHyhlfqVJX9ya99YwuithYYR61dTAOsfcl0IKIBF
j0Wb1dOuUI7cYOdh0uIcF/xdk3YNro/0KIEaSd6TJV1+yT2E+GPcK/KUoQIpMH17waDUK7gVpjFD
EvfL1JzuYNWdOlH31aHdhi1MELfrO3GTafW78S1z2uJvsxK7KDc7OhthY34eef396DOnBqZ0VIfG
0zj69Yz1TvpB0SkcEBiPd0ezdi1raqHgfKV5JLyzF5/kub+eWj0Fr+0mb7FL3Jb5n2479E9Dp1Rs
TzT7OoW6PUgzqQvkLjAevyBK1MsPLdeGqCLmR6cEBkV5CSB3wUtF8b60YI+5ZFcYvsUAscR52TYU
IEWdUhLaK/pljDgO7QfYT/XZ1NRUA0YCEJYUsSLSv25wPp/id+StjlJxKVgSmGxXGa56F+J+obR0
DolWHabx23y3C9fJT5Lf2tyeGV6OvaBaSvCMEfEjnAMvKhLX/cvliqCzsqSF7QHSwXeCw6i+HCfT
Dkib6N8f7vKOt+3J8kvbKoJmkJF+/ZjPSWiX82wXT2pnp0LD5Vptmo+1Wo+88VGgkoln+ZyZHiCY
y2pqCEkSNrF1e2KwahQVcyhs1RyXBSB/YMawvNTIqgq2ey6jykBIKqPdDndv+HtlORSvl83kOZtJ
ZkhnvPI8C/0oV+FwU5NOKWw+MksLVhRNYvGNq/o0Pd9cEwxV2/lt5WBKBtgFwm2/dlC279Bbwh90
eoBTmokrFEwz3unY4XeP1WOgKCoRFNVVITTHjkHonlnsthWJaOL/RyRz2mW6uWpBBoQcBrGHxdie
0Ftb9datZWWdEGdOU2acqEmVECZLpEsbKPykQbSxPi+gvrhid/gsYI11r7GRrrQVMpRKNIjrkRiy
U5BBYUFj8sMJFbGEwrsd0SgDcquCESmF2wrZWVYkF0byggvBmUi/qfY+LK1grF+73hyBwCPtk6KQ
cEVYQiZJsrnOCzHag01sJdPlq3pXnyeurqUqcApfU/UdqoG0+74PatqlD+Txf0jDXyHWZWThdWvz
mBME5wIQ2GADDxJpGzYoJtU5iUliQtDIjjfp6AhgylnGUDuR1DCC1/JTkfLR4HvX+n/iYbPDNv0E
SO8QFYUAh5qRsOodkqsfyzOxpPV/0oPyno8tXAZN3HRzfApJ95Z5epIimiuyTtBFTzYNz0s1jXsD
t5/CudBSa8gb6kdVddsyijrxJGFkZ6+VH3sLkC/yym0yznSz8bpEDvqEH1AaoKidl83luXPUpJiV
v/Yk/84wDtGpcY1YGiQgYhQz+8nweeHBYuwmId87kqVsLwErXz3h2hvguWiSbWsdvG5MyGaBVQiB
46ZitAJEo02LB5n05a3MPszMhl96u/OqtiGtsbn5XkluGWOUb7hH3N6pb95VWAtwpXRZX1jy3wj8
1OYDWju/p+YlvtHDuW3r8XDokaUv7clB/EPOF/8b5IFXdJfiAaJRgsCxdnjx/LP15T6WqZbazUaJ
eqaf3MiMUyt5dq3GT9IrWCnGoav3dzt+2WplvXbORNNgv8jtW1vB3QM9iKq/c6tpLSTANdY5X40z
y06WdLKWg/SIC7MazoouoA49IRGYGhghZUHU0qSJgEDmQ60/0emt0oXwizAB/lICImVGvgmlYVSY
07T3DxZHBnNBqGhztIKV2JuryI+KydhjEV9Vabq22v2DsHnJB9WVxHCJwI2VQSwKPp5jmO0G4JoU
M3Tn/xzlw4mL7yOx84zlcoovZt3q5KHON6/XNnxlU9O6MrckPB1HHB7zB1oXrjSIvGitQYuj0JGB
KCdLqoCWE7eYXHudHDlpaYlBVJ7TzDuA/Xx7hhkO4vC3tyfpIBpKpUQQhVNkMjBWKQa3uDWXakDD
7xEAABxA4Ts9TElwvE7KEZtM/FrhjtIZyaNA/4rgzTnQiksipWb8gzCEzLNn7FzFIsfCdadqSQCq
Dxuc1Ax9ytmDLQD4FyeSSkGrpHy+shbE+oqbrn2F81aHPZN18tkXYbr8mIof0DeOteZ+3H6ETqV9
F1+f7yK7L2rmLtnIGAeO0PW+QShM4JpOAtwoMcHA5hWeEaDq6iab3bFSJ7Sniji99q7TpoK1KaLr
5mp2FDNquRRAS7Dc1/9HCaV/xJK9XQy+Jp//ZXwEEYXa820pWop5jnYISSP1oJVxIv3wR/Ne8N08
565/a7yiBCTypORj1faQw+DiHqBSTXkTNWpzTy8mnzWVTCNOKZ3f8w3fZe0ojGBbFIFsCiS1pvWw
g3CD38NQ2VcqGansVSNoJnsa6GrXLSsZtsDGvEgTBRyX9nrkbjhJ7ZORELtugmWDjG88/Fu1yUMK
icS2J0+oNPCivUq941PSc4HeAvXH1mCRQSHP9wC5VV2E+1HOaOwhSHGCDaacPUJdsnlhTz5Au7L5
nedNKWqoOLXaBPtdCUO/yaKORuqjAClBNYJyUghUOKs3qyyhyp5lAOf2qzkqHo580FH/XXlyU/Co
+vnsx8H1yPtpsPZ+qbsOhBWjHV5DUJmyrjIGp+5UfSWrmPGpLyTtqxhwWRh+RKMFH05wOfiT5S3J
015ZA75+Mt/sAYNB28zkQjsf4x4iDhERwMVKOTiMXaBZcPHxdmZ+c7//Y/ExulIi76ZTVcvhhtdv
vUmy0ZkHeFeE8iow7WPC1/y3k6lplAWYvkKGBqAIx2v9ClZ/0z/L5F3GYRdh/+4iRwJ+Tc3vVMOM
sIwqx+MptPWoIYJKQXKjTslj98mShC8eoCq22PNrtEcW1eNkmUGrEYFvCjnUoYv4zuhTirIVRMiT
BGpG9SXqfJVFB5c2PS8wB9tta03kymT0rgcjCRjScV0A7jv5Pw+idx2Aa+gj42S9DdKFwt1MDn3H
rFF7NMxfSRGQm7UQ0TD/aXVHHJg8UBUyeiyVOVC52YKLtZJTKwlMFqWG8OFDcr8a1i9pxf5Zhqnt
EGd/nL9sIMRc4KZCg6lyzxaUdtrBuSzhJ0h9cNEPwJiF5NJ8077aQC6TRmaFSD5od/38O/1p8Uqq
ZdKZyDEKkIn0dmG9rY4ufqIvfBzJs1sRq9xivJdzRvKFq1FKWcnc+D3GQUxRoCjNjLAelzYNqAsX
eeyVY8BijPjFyUdfUfq9eIbFCjRwnxQrnDZafsjd1i/kTRZgraoRRq8q2B6J68o0LWJq3jrZy707
btR5a+M23etMpJmAz5ej5VU3303mYrbOfyNgyh2upoDY/x5vMORNJMBizJ2QVS2fRO3bcnYJH0OD
8/8+iRB+0OL/rfIwEgkgb6KSL2QTg7ord3tCTjEYtTJIc8kbcgi7SSFOsh3uqHwB3A1qWsBlx815
rpLkMeo5DmAz0LoK8flVnF8rVA7hxa8wrMtQ8DI1HubXzxxyFhP1cRLvk1ABa6KPC24ciL3/1vSo
vIdTtZHx6AGiAoIm5NrFW38lJRB59y++TuQMtSwsBiGoA78cjW4o5IMWcvGPqGFkNP4QSw/kLn0u
FoEpkU71r9tpAyqjk0seN8k72pbCqt4TcfSZp8Mcf7ly6bbXi/FlHbvfnThF92w0lFaB+wOzOoEc
B6kjrMsHEbCKFvw4sDsdZPwDnz8hs/nIwSBEKznVvUt1Z21TD2gUmv3XtpmRMMx0Xl11mk3fSVz3
4l/D2mGth7COxIz7EOPWq5wTfXpAL1EtQ6kS70rv13oTDkVMHigqfYWhpk0Q0CzSRhSjDNOEbweL
nISGvzDDhqfiwxoolE2mpr7I2JBGg+9JJuv0xXAb94Gzg/sGH8Pl1mwki1NoNS4OO98JCJtKTSlo
+VUDsW8UH4n2PcV4D+6brRZ0t8HNHm6CPo55e/YhTJ6b+nURGCAUIxr3LptT4LnSqNBXyq9z3X9Z
DLTLEp4gxzVkP3LhYETFzyqXsZ84GH8BZOEZsV+9L6R7frKqVBxbyBDA+rLH8bNAX0b9sWs10hnx
LUfxoUw3HV2RIwkfNXXKSzEK3GIsobiyBXgEgQHZGVdbVsaqy66IDR23igY3NU1ahXnQKxDH02e3
Y547v8fyMW80nsgBjw2O/1bUI5VmC71Y8DjQM+pGdCoQeA/1MaXjCjAweuBjZtnF+rx+v73PAl3T
gV4+S/D2E/82BnH1SKfIIKrTTkFneZlYZXIeC1vP9sxTA0IULox3cpTydTR02MDwZ/UlMKfHEN13
QU/Cdo1zJSzCwqkEFokedrs802hx1esZpATlVrwpkZKc9UyqcvEDWbMYbarYHrHOwFJ768TIPxmS
0Rz34fdpGmHlRe/KfPOAjeEwCtibK66lh4lFr4gT/CpP6sz8Nr03XfVH7/rdtIg0ki9tWumGrFpg
AIxQUmV6EmKHL7U8KfrgIvGWjUFOySdQnoDfGiDxIDKkwzI/YOpNf8NmOFRuXqgYgPvZwB/VQF2Z
WrJxRlDQEWwSMvGgKqCX29VyWtK2dNUsjZxD9Zi/vujv5G14wN6kCZtLtr23+/Rw2LHh2oid+sau
GHVkR4v4fDVxYVHhyMPxBI352/K5maJTdafNahlprfVXApbfetAgxQtegP7JHEOGiBfR77YTFkF0
N3iYouBv0OXcCTWkQPKyIFXgaTDdzs0nqMCOX0BAt7KP5StTsOEu1yyzwB44SMiBf/oBxmyWYloM
SisFjwZNR3NqNgqlMn9w4EHxJiccFraVgL4ji9Ztbv3PRsSSdOQ7LpIxtRoC6nXVKFlLpK6al5En
rF3QXwy8+FFL1OqJLYNydpXmZrsvctESisEqwocPt4BXKgmSh2LKf75OTOgr4bzBJqUDwORZVo/Q
vPC6VXuXnIXI2owO8VzdMM0Ca4FLPkcLEoYC5EH5RUuvyt6arCUI3N0wXgrOoegybfYOMhE0wafk
obEzujBu+AiLGdlIWkHUtZQmxhE6UmksKcRkPhhh58StDObO/r3opBLwSFo3nDPMqNn1nFfMAqbb
+F7dL3Vx/DGrEizZJEvvX2nQ5PDdMIKPMeCst1NIH33sNtMhDfo/qT7THZtZ6/5QFXfCpJi3Oo95
mpxXPT18fkPG8dQDg4Rdd/6qmSnTAVDTa6FyZAFpGhs6rE3nPIkj3iWBmXzkdvHsXWakz87ybNRp
9/kL3jgSyf6Mr1MWklLx1Qq+GCAiWGapQ08R1Ijnl2oh2k1RcaXKUJj+ZoL5FrpAb3kSVvhSr4ta
LTWrBxJOhlYsZ7BusIMqM+vsMHzt9LTQUpA84FAMl+r+ZJIfyrdlrMLgihq/fj9gwq4GGKfpuMy5
AaCQVytnqTboXKEo4QFTz/fhs5Ew3lazxmvVDwIbQL6V5Zh72QGUM0jqaMRhdkpNBIi0LPxvExu0
am/VR85SrMEHPOji8Wwkg/L88K71VBFJ+GiYRKhVJaUE9Um5MeWZ1QhLY0kV/PC1Apx2tBjqaIn9
1dFaOPbV2OZNPvVuLdtWTlwwuqrngr/HwDIgjBDJbIcSJfDeeH2uyjnyHiQfyyYKPBa3adoeQOvo
6P5UIL99xAuq9o6CY3S0FjorHc0WgWkflO+HCFp6XzIoWx5oolvTevYOTBMRHpQDfIJPBNx6cSOB
Sb2KSQDTxplgRxzkAGG/ZQ+SjAdnDib4XbcobjbABvRUlJd/ne72B8RzPvXGSCHEAKjjjMnp04mL
ODwPYWGPXOpSuauwcwYtS2E/qhrWiJEoEuPUkJqLlPpbFO3DnQR4gZyBAgtWZWjg3YgVZmnp8hnK
uOTMmk5Gz/MQUh4DtvqVB1sjvwFnsSrFSVT7R7FZy3/vNisGy0pP55KbAXli7tY4ueLSk3XSKj3c
Xi7TmAg6xRcv9+qoaXufkyKNqcGlndEeSNkWvdLpUNjuyhhzv0EXmvFM+Vq79UTA7+7FG4ZV3NlV
KPzcsTTDMF+6O9GUSfwynynYDiZmolJYT8vcABgN/MyMlFKVKk/PoGrvXuQhdeaVT+3JCIM0e6YI
I/MLZqfhJmvmZt5CA8euE91mMUDAXr6nL6h0OIM7G3XKk5avYI2RX7xu7vbtDxKNOrEupaChWPDB
aJ6pwVZWcrOswJrMQh1Mzeg0oulAbGev1C0hehDrOQKi3oFwYNPG5nN+IKwkdD2M6oBA91bfEehS
YBORswcPtt3GnSesgkFD5gd7F+IrEAjQu2k9Tl6uGGfs1YvMdWuqZFTeKadgsZcx2sOVy6Es7wp0
PQnOCnbVFQXIqIxU/2BxiS1bQxEPtrruP+FsvAu659fg+J6XMO4GlDlSgmKnJcj7XSDCgBF4bMIh
ZwD3IPsHI6k5gMPh4wnQmrfInWuCnf6tuJ9PJx3HDDjiFi2zkOCLAyW1gVXeeTAs/kIYEUjPrzHn
fELjaPrkhplYlua9VfZ4eTIOKxhamWVWIrffPPZt3Dsrb4Q5LwszhRNnmCHTStBFFwCXlHo/TkJX
Dm5uHQc4mRILEHrfZiWlRHPqCu2yIhI0R/2C1N4O66diV45Wojd76tHFHcb73PsdSY7hoXGylI+k
tJmGasym18evQbBspQzXzozUJE35A3WlfWjpmDXtENvQJnlP8uqFmpwhEbs9KtDhCkHdl5qOvVDC
/KxMmsqvcQabrxYcSjsG/ueoPIMjEQB8N/EnQ5y77sx1giJIPmt6XyQ9jaLnWV16/Aum7BhHwFAh
zfLbqmzBLBI046ZPGTNiPQQIHK5YoL1o7GXHHWwO6hRLtwaypYea8DzKbmaB8wmR6dFlZCa04MCS
Mr1UZv1lGaPTfGE0D/ZuqfMikPJi6hXW6I47oxfjauof6qK5yFgATVmzw4OMVePlFYrW1NAIE+We
6dK1cFGZ3onDLBbYD0lA85IbhHMg+qqt1iyRAJ5Zp6vA4V+hzfgVG0cFwz5/NMDf/64rpMV17bMz
AJultFaeydFh/pnWZMA7A1dav838rD4eUjv/fwAPXZr8hYgoAueGGfPi6CvbSG8sFDT1DxczERak
q0BofQPh4MeAbHpt7+1fkMxiHBC+zLfthe5B9OU8R8jursLPDtbd7Y9XSjGrF2qt/0FwVUqAiFfV
/dcz+cD4oZcf2/VXHGRjNXwAhLt5cj6QP8zxDqQGJJkLq63cvDDKIGWrDy5WEekVnc5u4AKsMs5v
23CnIs4P+vaqHMpomAx5U3964HAFkJ0BlNELPcQCsHq+57+Qx6vy9eIPRoA5H8eWtzzEuukR5+k6
BtPhh4d4ra760GBLgGsBHD7WcE3hLKObfckrDLY7kxCK7RrTTs7+jU4+QRNoQVRFmMlv31/cui8B
/JotvK9cbJLloepjmnBx0etvybVLDAv7C65Kh/fW7SniXYjGlvsYHyS9fS54OE5zzAKF/M9iSrEm
XvyhR64Ez9+iCJ8Ytn86WegQJvZGq5zL2wYpXyitlhROEzjBqffNB9UGvXqy/6htUHDNP4Jk66kS
0uAVBX+QgaCc+zJ1W3kiOLSRJs7n8Q1PO9hdZk+X/CMVV6N2UtUXunPwplriIAKwn3TUTktpD11D
h0b+BE8BE9XQtePCCOG8NPCJRji1cOIcQvmuQY9evPkTxQxh6Lzk8LGWvuZnsCkWx+E/cvd89otn
tn7KNRJmZaHqENGC80rmKgcTrgRIWoQKkXV1jUePdeRXcBNsdn7HlEay1cnzATapWrm+BBNFLIvD
MhsB8Q2XwefDiBP0TEAXx9mPuDUi2B6tHNHfRYfXB2djKJSkdQuuNYfBD8mspYJ0YxR9KreLJK9j
m/91kIOBHEXg9916fJEr0AFYw1kTRJZphKN1LI1GpE7jkTdjHmsQvaNDc4ruvTVFDmrBu3Lz9Pm+
M9BZPjKH0abmqy+09gWx8hN70wn6/XpCEJf1+vvgdUAPSkkHv5VASnoUKek76naAnC/lQ/7ZfIx5
FF0ifF1yujjz8r5d/GqMdK46z45jAmW7j5mVSBs7xO7iqNDzkK2JjYP4tCr73C8qQcYINqR2GYuV
QGstrivOVTCJ/XUCRKCYlS1ySslIxjpLd1bGHqxjhI3T+YEA85Anx/bkfln473HCnzy9KCfQAP6n
H7U4NbUDuW3p237f8q4GEHAPRdH9SWsxJ4svVIGNkoCkN5mVAcsS69lxxkwuUFxmTskPQdf+ymSg
r9NlO3KgXxYJHaBxlI3z8KalV4LPPC2nakGv1BvjI+y6LKBPm4r9PXKotbq0YfBuIF5ikSjxiqlX
PWeCiru47vgEZW7P8ydvjesi2hoYmodEucVsvmItgiKiyCRjq6JvyIK4lULBFBuptBD1AffyU+Dg
Y+EJFVVJ6qWdtoM0no6HiFZu7oxP8QJk0Xwx//+gOdk98KItRPT8rC8t9cHoMjLql6Js9IBVqboA
tPJR4KSLMw9PLgtjWDEFVoI6d0lGoJ/GU2Vg98htAlJ1sQXHVgoGReSL2ihsSagoPntGMqMBzO5C
yBS9mjwFo2wKBrcRdjq5L8jzs73WXVPS3olYdCp+eVJzo+Rr6tvCFPmCVJDfqbhex5YLcYeuAXaQ
fivJoZmvI3sjUUUTaR0fef8z2I9k7kvzkv8HxuH1Bmgk+5kHUrt7pf5LKpEaOCzMBDvPC2TYAK/W
jUhigvvTdxvHUbN8STLawKnMJol34bG2VESl/lHy2vjFxlJPdbfEpzFz1vXUTIPvz+2oEuEQppgJ
oZLbjuInUNWGituXy2jOpED3n2Oh85tBDwjN2mIVm9HiOjjBmbHtzDTdhsIU5vXrjY0EHP+6mywz
5R2fLrPIKhDv046uJ9YHwwzjZjrCMxmiCvdgQcUyCxW1qcnuH3103wjC+KcM72HKi6xyg5h+AFsl
vl1XrWgYrAT1WNerqexoJEPzE56vy0EOQgtPcFFTeYxbwFXs+uw2g+VrYBa139o8+mrzu79oyO3n
SBCksR0kGkiZTCjm9/xRKtptQYvEn62YclNKirrOJRmpWvksuJjZA1NILNonmQ0Dg/v684zqBQys
Wa8UW0U8y/8SHx2Q/pjXZueKyw584bmBz7Fyp6XZVOmnvyV/vXIdx0wSbzW1L3DoykzG7Cmo5d5z
tH+MWtLpS+qlB4Cn2tmDTz+MU/+DXbnj5C8XKYsfpXu0lH153DdSWumT6T+mKzP21gXJoeiD3JfH
rpCTk6ZbGogfNWXugfh5MgGdESKXWhoeqmhguDVOH4MgVFOJB1Lw64KrG1mS6iLsYfoE24c7Rpdx
i01lLncmH8yMq0EiuVMZ7KGHcDeOSptOjpKw7h7dPYdVxkPVZe64kyDhtB0+WWdvvduWtXFw7wvZ
VtEEhy3ASiHJuMN0EoYNwPfOECOuSq4vBbdX9ZZaYIrf6BslVUREU0uM50n8CoI1neLFhucHPS9G
I8j6ih2K/5OK9mZhGbF+YQyMoQKRLvwFvME3lts22UskeijrGErAkAVn9K1WT7QjASIMKnV+tRMO
lYNGPzDdnrwNLydXSe3tHbycoqjU8nMYJAwFoEpKbVN/Ctkd92qbQ9KF4epELEQ32uP3iEKRKymy
9Ff0aVSFNYpa0V4aimbzyVMbcx9raH1axUWkvxG75Ug6zSYzikE3Wwdt1e3LJQT6Ioa6K0E2ASce
1BfSgYDysYP+/4loAP2rGOIVv+/NGVRvvR0tASFy2KlyXGcMfYR+Ohbv4Ph/+BH/JLY+31EVoDSJ
V6AGwN68m+8tApH+w6CHUOFYQxfYsakKAiVOtFpSWVGQBL4sauKRhSGBigbp7bCQ8ze3gCQObmAd
Jv/i8y34dSYk+sSyXf0Xl0wpYkHls/UqHtjZ91/1edQRYxweWC7C10Dt8SssiT1+r1RQVKa3Iurf
KwpnIYOZIB8Qizcj2Goe2JLUUbtGSFu1FewwdQhOspM1e1iT7BwkePe6x/d6mSCyp61+GqOS8OwC
s7nS8WlszLR4kC+rrQclfsx+vrY9BF/NfYwk8f4koYulRk5AT+aVG08z0daP2yDEzUxJC/srpPKv
Fwe4GZqXwEEGHhL5Yv0fxkBYrE7Rw6h0x6CdU98DaZLXrXaWZs3Iyh5vgizxL/37Z3xMTfmc2Euq
SUsuVFWwqEgeZDRWnbENsxmRZGNfgft5HP65X4ChmhgXtiOhWbX1WgTvkdt4NeXhJsK0M/R89+rO
84M4ICmyipZIg0JtmlMBX6/jWda7hpHlItMyxBbzkgnw5UonOhYUyefPbM0cQkaFFvu3Q7xoedkE
/+Pr38HSHQhvjOAMQzAKBH6C5fppe+3oeCgPKj1QG62xaLfIYbPSsysi3Pux011RgZYRWnCbbKhC
KNZJAK1HTf88v40hezCL06/m+1xq277ZiM0LDkZ1zO2AMgvYe9Cz7qK65VKX50Cfq2pdX3b6+L4r
CZ2Y57VRVDFMOgp32PzxGvfZIyONyi6dEtYANXVXjRPWXtqK/34hw5CiQ4AMQeYBY9TCL/XgUVn6
VohS+NpTnT2yZiPTc1GxEUqHsMjgAtq3nCl13/QxhxMzmdvmRgYpwbZFXatsgRdeACBFbMlmyz+E
eX0JYGT8CI7BUnWPGDsL+dgacUHtevPAwfcuGnriI7Wm0zDY3Gnx29RmO6srBpCAqqhtTMFv+iii
dv+j/6a9t1vlt0XrdZF/xVWHnzX7Ui+Na+MNFiP2h6M6DcdfrsCC7IlWHDxm/HPEuGSpjYH45dY5
uco58UAPKsfdd2VoJYSF84NbLAyepuryNQS8ezDIYQbDikqq7/zg0x4R0jH/PKyZf6gnColginAz
hjO4+13PDXxGhYj2fg4vnXjGyeack1oDrPmePlH8q60GYnUeobKJO6xzGMUcDdZ9iGSn0EMcQ0BE
WapNQB5r13acxRZuaY3OlYmdyJTQbWTc1W2hnbf2LBjQt/sw0S2Ias6pvrZzLsoIIrSpHX+GZVIN
dNpj+F2+6chSXxiYdx0Rbntvc92bxJ4O2Nz3EPRDpzUw1zJAFcRtFknAPmWD8GN7HYynpN95r0SG
Xo6ben41OlwanFZ2a4gUuiW/j0l43Ku07C620lQ57Rz13TIU+cuLFcSYMOroFehoxxyk31306Wav
kpIG9+0Tdy3T4GfU5BKVLcF6pnsm2cN35h+RxzfmLCAwOu5vIxUfBeZzl4AenSYkGKd5UlE6hEJm
wcucuBuCEW32CIjLOEgpK9zchuUWMFaDI6vRTwyUM9SlJdTe5e3/E7IrmT6d1T6ajKTUA2nRmJtk
O83XVT4aLyVvc52iU8sWT5hlFayuaZEceGd80JEiZ9aV8/+L0uqMB7WrZktHgoO6YvYIHIiStfbg
auunMLD8n6nTgv4BqwYggddq5hV5kBjd+O04Op5S5w2D4Szi+oabBpLBcX93mhcQt51wYkyHp9Mo
l2kR0w7Cq5MGqSa4+GQME47GFXqhB6u9Fk3fZyLxzWtpcKjY2AMb23tYT1H2IJ01gxPCa/V6Ld3m
KMOX2EAa/QtXRVCFY0qLOUDIpEAfnFQbmle/IwgA34cYG/q8nPsKpOJDYUGxmNMPtmB/1vTVCtER
26wmahHiddC42C7+cMPuMtk8pQkMz1XbRyKbZJiMUFzFosNktiHJ3sI/uomppWZQaD3zzvvnWzs5
T+WLb98Ycbyo16sDT8NkyrH8AHdCvIhROFxuW+89vrG0DVix4mXeaz0QS7mWK5gYPw8H7K/zXuBI
SLA6ezNxxPXNh1BzMhDEy9KMeY4Aat4tp3Dxh+o7qj74c+oDdZw6lE8wDGbwrrwSFh7b0rJH3AJe
kCavx0NSNgMQWNnPHmeFD4dCAZt3V3CSVk667Y9/If/AdqbWMmZ56i/unFX9OSNx+OuIQggalUsF
5UWL8GGZFXvK54x4WLspboSTu2cAo5RFwF8N7A6SmJG4rCrHO+a330TdgJpRBM4GEgR5sflYK6Ay
NvGR0G/VOXtaGLJhBPT0Hka3gb4YvceR9DcgxAPUNbKNM+KHviFd7mm56BYtAXuR2q5X1QfErkWE
bnd1dWJR4rNKHQdSQA6fWqGxzXEuIjO5P79jb1xwpZB07vRgHvvkhPLk/KCX0cCzJcBo1D1Qc5je
CVRqfSCYWJGp21IgE09oxZdwFFLxPPwO+iqAwEJEsFIzp+DjXv/Q9GgigP9hpE+669x6p6LJWVIy
dCQY7dGxcGPsZcpHpgXMQID/Fcddcr6jqbV4FlueX1QOeQVNZBvQdB0bi0HLMfpx2Mob+2njuZ6Z
By9alX+3x6Qs/ekVtZrn7L80HDUvNqfpbALvI/ZRorB8fGuRr2xLyXGIRnkCTzCT1ROA2P04M7uz
MxkyzUxY/KiViJLF29M2PO32DG9ekugkb1jjbJ7VwC24veisFJpCwn4kkM0Ux/HIwbPbpm4h/OWj
amjajj0iwJyAi/Tr91909BYc+SvgIlHSP9MHRojXRtsrLIcWcNRK1ekSeBn2nr2o7vaeJQaInGrv
onv5wgcPYMbSi+7vvKFeqJQ5Uz+HvnJRfLqg64wkRUxilwSnFQMpaVXXJ0pCm0YbT55zP+5n9tN3
MGgFXw5s+OnZTBLB9k98/g8Yb/5nz5Kc5mwOWHRp3RmXdzasIB79JG+bEV8pPd2l0aQ+agyjp4vZ
BzcW0kOOZVG49vyQD7/K0en1yuOD9kH/p17vGoFNZE/gz1/GUNxU3tUgDZLcHZmctIzs0+USaC/J
SMEJ/lI9y1t6LpHAnNuCCld+Hanl3NXjg7ARWDwl/ZIaPkR82jWQtYvwskEEsX5lGqZHRo/5kFKx
TVtygfYDHVGTypA69gibntEfAo7i05bdNyPL3y7pIu+Y5ob00FVYB/7xOu8zW28xcSt1aizTk64I
uBFGiTBYbp2Ns/d/+R8kPnNa+zeJwLweUYswa9GyaQMEVSr3Nup7kOLRB2DCNEzp/5uC5anwovHi
NsEcuU966GfalFXLhWVjuNgjON6gr2BPLeo6RiZVUXduqR1+EGail55LRfOGCUaFQW/wyLWBmC0Z
XlePQvo9yTYCASaNUs8q6gwrrfM5koGH57Se90PnVnhMR3KGCtPYOC9OpruoIxHDP/wwP8cHB7Rd
guRv5HMefuCiBV5LQWM0xJvcqsAI2rPkNuIHfa54stq9Kjl1VH6u2oSsTC2ymdhH9V9nJJNDMTOm
9F11AhtD+sQxfDHUb4k58uL6nUbLJdwHcbIqrhhhtKjh2ABuzRWBAsOlfGGnq4681SY2fuAMYD42
tt9X8bdYaVj6QtKhraKg1OM1/Wo7zWcr1K3oWgUSLRx9gl9H3hbEDSpji+e1TDGwTnxOZdYWm6/X
EsOvSndkfDGHFEUSMJJobUdwilkUWPejPPq7WKRXhyHbXyynQd6VPnlJtXVSuLiD+do2H164zL+j
uQUuavXfw8Bo4bde61elXGw250kEQ/jgWZ0iLA3m8g4fe16y55N/1aZPNM55GhXjnHVmtvFkEOe4
kL+mOnRVbtoZDaXeKPtuVKIXXm0OHjtdHyiP8va8ZdXec5hbQDvUDzdpEseDk8+EneT8yUfuHUtk
yiXViDsEg0g6C4h7cyU/bVn04m8KcGBdib8qu1S3WlcTts/StIoJFNq7Qcqnvef4vTKq66ExOuhS
eKr7wI15fH3o8dwLiBr6Q3D3XDbkuXDY0NcD2CFaXgLd/BfDSdve0MYtRytraaDbtfrNGqThDunb
X3uHZk5r0aQgAYg3UEu6RFloN1zCHr0onjwMNGn29npjHuZ6hQ8BUl9mnLu3x/9GQ/CdwNYrc5kO
qM1z7J8VhWSbdbienCiedJnpC0aJvXIrVgEovROXyHKNmTbXpx/Mm9nanqiL0YQ0tNWj9SGPsjUf
yDzFbcyS2lOwE85+gpQTHbbkjzg6sLGZ96iYv36WOw6jbro5m+cRimAVpDv1Y5ZPr+UXnnMfcNWq
vI5d3fDRUebJESXdWp59xAJMQ1XFOx0yDzsNw3D3f8qsM+k1aT1WySoe26icCQRMqVqzx1nDLeoT
4z7rg0flJpPkRy3MGaiij/6caxb1KTS8n3QSbIiA0n7VIaRsbgQZHKEe5CjP7yNQP2xjlnYjAbGH
iTFpums4tYAn94NKVZWPWw9t6VXj/krxoXIoso2HzVhHf+5QYjF9QcnxUEXMBmf3hf9NwMoMTNR4
x1YuWtMn3a6FE3tPQlFtB+nHhaNNnvLQvNju+IWT5Ixxf0hLaKKzGpbckv8k3xkFsFby9zBwMQqS
0Eu4aCi1Ol3zlXufe6QPeTr2H4nMZecJaDaW0vmdY4FYLCmciNtl1WfU7Qikd2HiSdRTToCNB11N
ABszTRuihepsx45yzMD6weNgdo3A8jU6xW3VGnzjHCTOwxVgd4Vr7W6lmtrKj6aFzfWQHF0g1KCw
pcRkoJ/dzf6fSJUL5uaTWr32tapWiF5DAocAri6or0pMrEpiZOlw2/6Zmc7bDE9Mp4MRRSl60xqS
qGQmBLH+YvZi1mnCMXoS4r8Nuo3kYrogKHi+lwWv2SG5Qdnu5cvLsGQzi9tzz21lc/E3JdTr7s+n
3edk0TFWso6owaXEGsgnkvGsR26/kDbKWqBlAFhjWmsb1fuxsNOQJzz6MEzYMGnZ9H8Ye8YnM6si
yVWEjhsoJUrUJpu4vKMxVsuVKCX27lGryGG2B8/aPWhB5Lx0pfrWg2vp0ww56AGopikIp/fM+AFt
ZpRxU4OFOOaY7vVgsCRQlHG0w5R1pbeB/Atsv1ftlTm8ZCj1HP9OYm3foFG0jkyFAb2mYX6sLxF8
yB3hSovS0MUkQ9ujs9vz98n40AkFzjSd6wbJDF2GvhCh666G893Mv2gTZdi05bAgQTjLDSBl1I31
tlhlSZpdL6Qb++DGKyM0hasIuUesP3KXz7T//VFFlCLNNvmFPgjBf9XYM5hGXICMV+ZNyxEXUR0s
ATkw2Xeg9qr7zbjnA8yFAiXzoz+QxJUac7h7GpfhLTBDSAb3CUoemOL3pOcwN1oe+LwIxK9Za8VW
s+UAhvwQs7pXa2w1chpalMV7fW5qU7KvmxjzCr8G3hyhIvoaVMen0x1/XcysEJzNbLInBN8JkPE/
UAxcg1Y94IUl79gjNk1CpoDdfo/ATT7Yqg0Axh3Z0NNiO/o6gQ9bfkjq83uzBlFozlmB7f4HYwh7
KZOhq5Ek+vDwfC5NavbwJrotWc8C6ZeqolKA1vYHbfG1ciUb3g0x8YgMb78duNPT5EWyUbn5xLEv
fLujoV9F3AMXf/DuFsQq8CtNPFzbGsd6U18NNfzFmjPxdNRYlORVg5TnUdERUcEc3dHNlonYOAVY
fAi5yqTkzJvZ+VTe0x+gdmMhTIt9s3v5589Hjufzpco2aJIzVisP4lMRVd0zvfkOk0OXFsX5jhtK
W4iwAlhDI7UpXBmH9jR1l3U/Wn6RYtlOAv9igX+p3Ci+iIW4ptUxUH+mk9YvsMYKEw/xUxsxJ9/A
p7WMxa2ZnDMiVxrwSYv5Upj8zFuPxKyskndImbYvIMXIKR42mf6AMtscHjcLzBwa9Vfm+kpw21dI
0pe7DaqZqmRI9Jg+2pi69l1PipX9125Dcj4WBHdVlbpIZXox0K3/2EALjrU+vK4yJQdZZlvXRKZy
GHF4p3pynt9ONJQ2D2OgIXRZoV4bb2PdZf3Azb6jiJu+CWtC6IZtWE5/j2do0S9FN4WtYvhvZCie
WfGmwCpv0VOMGPapS5II2J1bkoMC1v08zHe9N6PgzrkIlGxfcNk4zrDecgDg1NY13wfgLU1+WtJr
g9XuGV13hJWLH9Jn+vtuCYyjYtfCg2TkorBXI5SC8Hy5vjH3XZscvXTvO1s0aF3Y6WRRZbzKa4YW
ykiQiW1BQ7+EkAUZfd5xCKQ/3mizhW2gYGlV3WQJfP8W29AThczMJqNQqShtfzRxiiMtBE/IpAdP
TkB4d/1PDQ2rW5HeX5oZbkIzOwauIsaEtPSUtxE8v/6hHz1kzX4vkcrPvsIK93FNGQUCPsXsIiMp
EI2PcdBcQjkONBZ6fpaY8nKp5Wy4FXZNd+7g0FetqS1KBe8X5hrYsRH3rF4notrRLouSXq+EaKzs
GUkFv8ckzrxxOphgVW9ILuABoaJVm0V22lHRo7CtalWXQZXR7uRL2If6L1ttLAtkpmDIHiXao6zL
oKwi2DndTq6xn/kDjshg08rBQmnaVB4eTN9ivuJTktj+bXD5bTwAkKwr7yNKWhjd2V9RS5x1h7vY
PfvvEdOQKTTzrTPWnPzRXri3UhCpryVomh5KTWJ+gwE206NAQLoR7UMJOeKRQtwxCxnnWcsP4mlv
ufSCAtu4p/4zVyT2na5JGBDzmJXgGq9TjkUAL4uJCYyOlncWBfa0dyHh50Nj5O0dFvuWn7/4asKr
307afzhUusqaliTegYVbtye/tIa14Ha2j1PJyypNu+XGvge8zjZdwZOQbB1jDOAV9DOK/R+AvLUb
KVEAYWbcmLXfQl8uaAoWE9hAts9mqCF4iBeL8kZMdXfPBQjfbG8Bw7pg5nHpEyGZE1cEAxktmzbB
hDQeK1PQKFAh0EBbs7s9BhrWQh6XzkQ3RbvD/SXxqQQdDnTr9idZ8a4+AmwAfxBYPAz5urJTbRY7
Khew9Yog7hF4GKPsjuXnvZ0OsQOTCbwwwVZ5sMs1VoPFcG+o8WUol9nHdsGcMtTphHDaZt8Ah4Z0
qCbCLUIkRIYC4Ll7lkvMwZwSZxXS3VDTBVgOQj3GJN8R+alUIQJZWIXae/dJ8gLgvZrj6GEL5C5U
ilSZTsBxfQUbVEKQ2Tx5Jrh9OgwKjrkDMJcocHb7xzNH/OMXc9ChPJNDh0uzmlwA7zeAfDtiR7HN
2j1GMPYzNSjcuNAI0ivMwlIhvOw0hkl5z6r8bI7lC9FT9wUrCvupLO/eYnaFiOppaXdknd0JwDab
67rs7VKzY4Bj+iP7+Bhd3UQ/zfViK0ArQBxHsP18D7c6AMcl7xfFMRAI5FjZBdGSCjvaqtmxU8jJ
3dIpFPrgDzdDgRfYUjfE6cxUpm5BqGuWiiPDGhD/mK6WKoSJTafsoDT7jKaPrXXhAR++jgHZ3jHt
NGbK2LgsXj2h0tiGm0AK902F+t9HlGXbRWYmOMt36d4YEUfvlUFNfGiU507oIifZGvsw7/d+/ttR
Nt8N3o+p+kSxF3wWHp7NTIGKMFyx+cNw6bm5x+JrMJwMF0ptKy+1YNSj8jurHZfpuapFnIRh0jLM
5GVc30VvnTV0DD8TyxkHJOGV9pZ1LOoCg19oMOYACeT592WDmXHUcVdMpzJKMsWdxGcGhtcTFO1c
gSdu7K2fTRiSTW+rxppiFHj+sI0vK6ehF+vmd6ceyeuLQo1w7RYXt5OQgMzT2RIlIU1nTLTw/JSn
HRiCeSM3/BWVdJ5GJe/mFggpXdjXysxTtYfFl02DE0ndy7+M5v290as31t+F+UMt+mtzEaroJJ74
kC6ujsVATH6cNq90BXs8t0qF5JgoS8iVEClwBXja04R/Xtz685yWjZ4Lz9XS9tMvQtG0bjV0njBF
nIucK7w5P/iTIw3RMQiI5aoOoe4IBPgUj5xW77OQVZerYMvRGE1KvhX+X64WQboKuyrt5rSvneZ2
A2MQJCskrC9WwdlKLfC0n6wrSEtqYvcitsr/G0LqfGhmMG2G+O+IJlo+LH8Fupj5Yf7Bt8UOPMcl
N34zF2DgKc3wpn6BQ15o2MIt+0yOLq/v+artkXIPBXpRStaRLM2Yz1zjpowj5O2b1nNBG4uGt7um
q0dlMM3hoJrR4WkShcsvU97bZjYBdvHRWX6D4VWQux4YlkDHSFq0BlnJqKGAQ1HRC98VzRl4TOa0
hpVkONtiiq7nNFSj9aPgJJLdSGXShQjUg4CKd/1rA/ZH2mUZ1bHG2YfjB2J6z9cuGBiAJ4P6xmgX
yo0H9CbKAWPLiP2bURQuUc9OKN+a5glz/YRpx2FPIF/QaCgM7rdnuQzq9862QAwpIIVkW50S5MCg
SW3Jha7EJUtRYYWhE00QW6PXRQeiNAvDFqyOcvnbCvoQWGBGeukXIwV4WYXl1QX7DZtqM9C/KKBJ
WzBmy5H+5cDNCsxaOc6X00MtgUmcNh4u2rd3ckZ3dU/JqmudNaPP6Bkl91ZIJJvikA77g9DzGsCP
VMdk5nSGqwUlOsAIHOJa6Lmpw5R6ht53hCjIs7LEIMrAezYxof0Mv6mosZ/kPUltGTJIZ6f+Cvnh
xer2hAWSsGfY4vw1VShcmTesaLCqVaoSsOb0DxJnpQDcBKkNFfD6JbZVh3qPRqsKi5HD3P9tFqr2
kQyuk4HiArXGG+0bqxkG5/xFQiITWhXOM1Fgq8fs+GGtq6WBKUaTtYKkl9Q/teZyDATwt/t2GQxs
0LBJSNi9K0xIm8v6BKJj9qHyARiuaFn7Di2c6ewXw7DzIKaEmSViAF5KtvrpAqLLP55efSY7ixPX
Jwz0bG6fL6T37GaMOUc0+MsMahkAjCDvcGYDjv/AalT9MFGv6u2ohi9HbMjX9tNq6bHUseEjDnbo
QK4PRB8Dvq/OPIwiG3Hh6ovCkkuZD7CDxBv7Hhfu35qAoSlQhHuXIYapmbbL16RXUyVd/JjhuEVD
KhPB0vwP0rcTF2Kgc5jCIqHPog07tRo1q5GyxAwTn20D6yDuA+By1UWZEckB89qQNYLT3UpJgqd8
gXImis2Bixc8M6W+r/TSaTF+pvZtq8du3l/ulLt6qVRL8p0SC3MVvlz+yAUWuJkJqMsfh0WWi5fP
zsaMu7y/u8jDatHbVUITzKrGNPqGXWRQulHyQL0gAWYNLu/hjVyyXvSRvgx9awrLPfGAGRSE95rj
fsOPQZhdjHAO4MweXlaDS0XfCtg0Di7UGd3St/5fO0GE0jqhhyV0+elJodkhlnZo69PE+x/+10tn
0AODJYNwPyAbBkgG2seC4Znv9P9rV2YwOyur+4ua6Ehal+uBv+ywNU6zuMGmbmOZ8TtTmbPmNAVw
xIo+xETV396TEg4MMFZ3vfZKYMkpmzLQKouW3FrD8P5vc/IK5337cfcEQzYsK0dRkFNrSh6vlmsv
SGccqUkuCx+LORBrXgKpVSdSGGbuz8L9h5vgAjUriGwWFUHarvngQjopty/PTM813Kb55utvPMGT
gVrQ9mfJheHaLmeVHxDumMH8ki1/znhLgqg1L1FEf5mU7znbG6YQ65+yFoflrIqkX9EFPrgA25wA
dG72oLACdp64vCWtQYURIND6JLMjl2Rl3NAyU7U3llQ58tT4RgxG9LZ0syFgn4vfww2wFhK1eUgK
aTclNvd76nqxd2oBM9atIkbWCS50wSkSWqoWJ3k8/RAv8AR2QCzoavZX2FxtaTs8OG8Nve6vXdMI
pJKlho9tb6ySL99mgDlDt3Yo9vv7jC2HbsAglEeOnj+5w62nd6Ae1aLJ8KHydl3O5LlD3lg7Tst6
1iykApmfRYwHFVl5/1yjORj5Ypo4yYbFws6k2ov1fC4F5FbQGP51VnfY4CrxrLr8vfmn25C/F+Oc
JQOq7Wwdmee5qinvmp6NBz77EtRNPC5F/ZXcj9CKILrQD4obCyEBkcPoXwO5mQ1UfuTo/hPZvyLG
IxHFeku1gaUIRFgmTYyOHb3yWyeMHxKd9x80ddbW5K0qDa0Rbu1tyAejyeaiPFwv5Ehd/6X3CcSL
6IvNBzZ2+W43UTDrmAlcplYZXP/M0xW6sPOXKSCUYCi4+EA9mPAK+GO+hXS2JXzFSg1pac6t/k8x
+LfgeyJzM1sQ569K7cC7sr1ffO5c7/XMg6zzIEPjRLNdooCa/BIoEzDk64peTAolkYvGfQmwdr4W
YfXzhd8x9nddcxXg6Qnej29cGSIfVq2z80fSRuFbCT+GVma7EnJsN7k+ysM8kOk3gmPPeGpEwyPF
Y7Sn2dzBPindwLG4r6D5B2GANVEjg5jymFS14KN189Anc34lZ7UhiE6A2V4RzaB4xOt1raMNlvOG
OFJ+3QSfDK6B8uitnAE8hyNoM8YH+z4+jomBH8kvSPGTUA1Nh5zLbh+Hq5yCYi1K1SXwKiaWxRvZ
FMN2lHQrQ8mao56B213TY8I3d3I/774KUCzKum0XP6o8wa6g3cci3bf1IHHYTr0HoK14e5bzc03X
cPvynmJvqBU159sQmyWy/5J6UGwAMaNYRfVL3A1BNeZncaOYejFWZLNtYyUK4svLvCBP1qWqflc7
CyzX3Q/TPjCEzHpm+ccNSW/WOvOp17p+N4BpcZ7F4tioa9peVSLUcJveDurAN1AIGGWnmFeAFN91
tNzYkfQsVW3or6Nh/SrJ63zc44MOl8bpHmDWE8evksdNXVJo0q+vnCNspBq4AT7TnGPYrIfqXIXn
gi/tbOIBw+ZfCF7B+X9S0cWRmXweIh+SaD3w65MI6mVQ3v0YRrXCk4+LzQY3YE1ZXJ85M4zUnknH
+UhKtL+bL5r11vKVMYL0pvSHgLNiORklxjnvxsO1PVJNo4IWAsLmZloRcvwtSqwUQbNVlSsA7EU0
PZnVkAFHE5dxcgMjT5muNICRRoN51XpOyGNtnVsQ9o1ij+MxDJqhl7Nd2UmjJJCzTmXYTjfURFn4
TiQSVxJa3D+ovTbbWldcVj9xpAyjCU4wQb+kzSqZ1vESZKcTk+qHM7eXm5Y2UNmbM8AwWL1cd8En
W3XEJNGW0NxpHK17Tphk8ZvemdS7JZGusZim4+5I5lWI7IMCjBNcriB3to4xC18ZQITWxyx84hMh
+sEEnEroxsu2WY3BDP+3oc0tqL0/KBJ5D1F+hSMFe+f3JW6CYqrFGPyzHHyI8uAzn+eU+W+ojvwc
twRXVYSQb+5QeAJkupa1dajP0zMlHSq5suGaYg/GTBKpYxgWPlzvGiIdNxXI2kZ7IAfNfyRvIY7W
DbzkbRwSiah9WFj4kSHZiXKIG9pxLcCwlYJZzHeQi4M1xFTp8K0cicRavT31y0MCH/zKwkHkqsR+
0aVyd1bXHuiJsiZA+GIrI1if5S5NySQtCZX/qvXIH11HQQ5IawBD9ulk4GCj0hM/kw0m7Cd0uDUs
YjGFhHy0NJe0YX9Flf/p/NnSyG4bn05cMKTi5zKOUjWstjEu1VqUY7/6GAokoZ5m1OB5vSQxR8fE
g0PgcJv6/8wa1CtRat3/ggdN+AIfpDFyBNM8k9JKr/oaobuoir62ofhYaQ+sv5NeW3T2JhSzzrxP
RXeAmaRvLj5sIJLpgFI3E+wHnIt7mSIP4JnNU7vbt/chlQP1YavoSWLKEU1fdpjlYYazlcLCpywU
barEgBrhbm8bUvGEzL+nKZ0+LGAfdB0pllKxuoAGa4mcDrleS/2ioy7gIcgj+EqUM9COlAwkfUzF
r/BWV7fj9YLKpCk8U7+wMN68YMSq3z3jKrN44aNwWr7bsKZwsSWFVrdkoQRFgfVU3tINn6kOFdFb
7VyHSFOyoRmGeEpgA1tc3bR0SKQTuUuYqHQhAbI78aozQGMmykRY6hqlxAYinzvvLYKHBgunvv0o
jxb5ygK3bkehJRWEzJA5hbmwG/qgKmv2ZoV8LeCU4tRSu+2JpIusuQvg71mZuG8/EvhyfNZBs6CD
ge6ygqqsg8sEEwuIgFlg3HQsLzxXOVP+0AXjVdyZZEpDmuOp8KnarEyyB0xY2fB9CrVXXrPn7ik/
dmn7KqUrP+2o1lyb+Cs/+6bcPd1E+9ewF/oamJCPl43ZnlIGOnb7qOL3f1OcWOQ6Q86V/cG0v91r
2I3yWj6bbPRlMIhCa+eKLHN74bTWBeGWSTyzeEjt2RjK9cHh0KSIFeZjNyTazj+f3V5HscNGUDwe
+mQSEsoKeAq+D1trw7YsQCaMWbryJg63ho4wV0u8eJOAFiKxbfyqGTvwSoZtl+XhBpQ9aPtwT+H9
+1QD5BMNMs+D/AgeBPhH3kbfYxrH1t5NGyh6ZQ3Feuz7Wsi8MX7ZZ43O1365hYjxzTekO/LVek8s
dK9KtBkSUVohEzVfEbrEyFH758WBM2eMfEzwNELoFx5c3gjIL7VWoTA96Xs0gHR8L+KyrxEjLZyn
0G6VOeIFgwzvkkHgEpkh9SbBLBoCpCwMKp05eXb4FDwxQL8NTGymtlc/iwWmDgZQIFyMVILZY+Gn
+Yas3lT3v7XlTVOi/fAcm3kFxQh1BkUxZUnzNoAY91GGB1HlXN0wT5WvQofsVw5BTNwya4giIo3L
yTALNGmPsWrjFfULZH2u28QuZDgv/pTxbApZ1ASqbWRnsr60MYJKXZk/Mb7a8wn7ICmPUOhXGeDN
KQzBa3Njuu1HUiZvln32x7KXkUyk7CV8dn0/sU1/oprGGL7tC2PUpzOjG8YoZL2+NtBCD9vRb1HB
IHWgritPBAB+fDJG6YhnB0Hj/+ES2W0K8BmfXiVCAtrX1EEtdfVblLvFx0YRzxxxVS+vXMefDZqL
jOhXvL2ScwV2cfDLf3qgOrl7Y9CbvOwo+6pm2Tabstyba9OgAlEUMvjm4j8HgG16qnBC+gRBKKOr
8rFqwbZxnYOYJIGtxQyno0MPCVWfNhsw7tgK+L7xVvMM1zu3moT/Pc7wRqIrjFDCO1hOtOuUqKeq
phUll5uiz3WBB0G3hNeNPzu3ML6FrdlIfLiohTbY8TZiEmbmpkfIrz7sJzR0pnjy1cpWRZyzpCtA
zUhu4yqygzGcNugGYwKkvJZvjupIb1aJXcsKjcrbZk/sb6x3R8sl0efyQIz0X4PoxjRVsszUsTCY
VHYTZKE2AI0ZWo0OFN7n42WTlFeZobvSqeKMjyJ0PgyL3XP92XWkTGZbeu2tstpwQneBXQ8Oow52
7tXTgwUzcW8ozi8oACvlUNZV/6oJrNtxtgmdYlc9E7phgc3I68ROczRywo/dUVEi54xUDSlHPg+z
9z8hR/sOCUdTk6JahfF5g4ayhHeglgIFvdggM1d6b962nRScQElugWYL3KYZrOMyAHcgtlj85Xy2
tlGxjvdR1XL4Ax8oSpwpU5SQKUn+Kv2lFZKmGVtpaaYFXKpnbRFdjzz08UYGeaZfnmKUoQzeedDK
WJct5KgHCw0743Um3Fn159xAHwxcDTHKqwHH18Z1+HSfrzRd28opGKOwOQV4Vg8oGoH1zN9GBSIZ
2S31hHCjcLgCiKI+TR4MQc6sLS9VXGeaSMlhSrfUyaT82zS7Bvgg9BBBXPICS74vIqVJXPAf68G+
U33xnnwQnS+z5iSqic+7TseEogUpYYtanpuwn0nchAdBdEyhXIiRnX6cjWR1R8cnSkfgc13zb3md
YyBUHpdefaFdA8VnGV1YeqNlQ9HTHZ9x1pKkiM16HzExldcObZgNImQdcQHxwke+OJigo12QdHMs
95ExILODjy/ehlLFi8umenrxKJTjUz5nzsLCI7Z5eqW3oEwVpbCY2ims0cdlsLzRMsyMTkeC3vXd
YPpiInJn+HX0faYfP4W4xnAx3K8Z3fgahlmVCciLNXgoSYD4H6jieDMB6xjhouAWEooP2NvHajsB
ZaHNzkGOr+QpHIMtMnYBnuXhOAIxI9zepfc0ata8Cb5r9ZcL3UbPBwB1nNU4Tlm3+OuCtTq2mbnt
ub374pW/p8JFdZ0MrmL/Y3c5hTM2Wu7LPxg6+XLhSvwwI76tk3l7E5AcHSt5JaK0nZKc3eBAmRE5
ArUcxV7p/6uTATgOAntCFlmeTB2Nb6PMrknxLuMAmJRUUlh2W+M5sz7h2pBJLoFpihC12OvWHkDF
wV7IgIFo6oUOOp0iMdxfIu5Hon+fZY2gXEnRTVyUnkIfamD3nWuRP0WDVmKufb0WWqmcfi6JukrB
4hBm6HISLDKLseTqe9XSdgtFJVcLfH9vpd2g8fiIDJy/bxdg7ZSBBRwdlYGN2FVFnopppeLF4xHo
2SmNxffCJXOkdAVi7yWRR6x4uFDTXtaM2bC66jS0xiYCpFwHNHBgjN9BUf8gUYBJ0MF0PN+6sk4+
JfqV5lYysLjg+ayfvOm967+YX+LxIYxPfY8N+NB8IUwtlndV5pByRZE8hkKjCCwyW+cMQDgxG56t
E6/UhGWqQhZixxyvYYK2ommEbQKwV/Q7CesYkXQfHVjtH01/QHLSO8Tek0FyQy7jDISZGCe39uTb
s1gudxLKsXosuiZPW/GnRdnIHFAl5ttnQRH2v7MaknMgbWe0H1w1qRYnQEz+bjG2kEJPj7IVjz0S
4UKJAgkfLBOHV0TOoOsOb0r8Wh1LI9w8XlD0zWN84sJlq+BYUoKP6FSt+pS9IvXj+2ExxTxyX7nd
ltREktYeE+jGTMttKoQMQCzMQ+e+aLn/0qK0nEtySkTJfA1XpCNLsJ+JgNJEg1dkAgQpzAAVWDTd
yjOTmXtCr2sCCt3GXH2iN+04bvat7Nsg/QkT7AixU/zI0DKnhEt0K/vL2MyOPuzoyv7fsbT2xAOc
vVzSwIKJnf/W9HAAWZRtNi0YosGz3FPQ2XXed5IZa1g6cj6AxUUe4pmJYMCjdeJ8nJtbehx1kHUr
L+6ZevDMLTxDE91oG7IJTGsCZ4vY2Yao7wz/fYCh0tJHm/g/1als8b58kyWUB8RfJAaHDqPBe4pD
8siNgRVKKv3/UukgsymWBdiVS24Y6vIFLnm5lDEmDrEenoScoUOTkswy9O3+PE2T/XYvUtiS4nhP
a2749XtWPDvSP++8K5mQ7YkKRWCbOOaqYyR4U6ksd+868G6w3ISDFdNGbw05PcHDksZPDLJQTJef
7THfo/F5eRwO2eimAOayKcotWO7VPEMMyoNaMfWk1QhCe2PTZJ45V9nc2nWWJLnNAGhmSFUWnb+E
m/zqDiaTPcdfvpYcBRQTk7ctTQR1wWpI1t2zYwAVCqp5/ROyUI06boWP2oljSKK4hg9+YWkDlBGL
rpAS+yJiqiQHm5TPCHO2WMDdR20IIZn1KgE4apMdOxrJ4aNZ6IQbgRTHMP7Uuax6FcCFitH+Mqj4
SdR1a47yuANWMKrdanqSiaYX2UhMrO9wm6JD759K//+Jd1r+xbLjr0XHMHKjnEx2YojWGagUUnJ3
IUmzftF2XgPdfVtuOFfE2eOAf6bzAS5XilgMFzBIljyPDGSRnB/mKmnD/aOdpLFJt5Bo7pMbNcoZ
rLAo72xBCKzu/XF+qOdnVTo+qGFIZoTFIIUJHu8ky+GRXOCNW3nOY4c1nUa5IMiEz1V0gvkggtgB
kbDBWh7Xe5cpGn1h0r/Yxzp2NEF1D4FTgsVSKc0eUs3PRPOmo1BAIukDOV9m3MRWAauVBcQZAvUY
NI+fiYgMG02KozLwF0uXwU6R9RvU6klonWmv0xTfS8iruFHtDhp0ZdW00i1Hvgtqy075YLlUwKzA
WK2AbtmncwVg+LNYSTxQRsqt0q48EjDg++9ZX4umj/enMMYtNu45E3RzeY/X3Kd5d05VRxBHbL0D
KBmdMYfreU18Vgpge35hRsk1d7rVtpr/iYbikVwoCbvmUNTtIBIUZmppcLXtQgG/Me2NmoHTXx3k
+xArRUkgSOpvzwhbda1SdlrOttMCgk+Q1F5LDD057UcjoMkmoXaGbLFDang3FmeUp9wR2FMVUxMa
As09QLjWjpYLl/jHrWwCKuCAwLTKizUkFTCQJKSZC1WoidZxKIkv3gNAIy2gXMiKoeFie6EE9Nl+
6U/U5Xrq05tw4oxFN/L2Uap9Mka6m/QVtyjhZlV/BQmwffiPFyiYsWwYvkkc1RobUkCVEXBw6JbF
Q9nsBfBVOM1ZKjMrYonQMy5MteJJW5v3f7lvSThNYKhoMy+t78ZO3PyDSDEYRA8dlXPmb15Zy0tM
U21bN6WAowTdhpJzuNoAU9Wf1+HLo+JILs8xCzqVktKlRGAc+U0sjY3AlkwCD+ixAKH06U9soHay
U4naNS/hKeiDrLxXqeeq1SRTj6Cy//uyk/g+5Ruwms7AXi8/RhahFgfYNE0Gvi1K6T1vDupXSupg
6sCNLo6FDYosL+9u/1jJyYh0J4KgV77c/w8cV8u3rb6Je/tEsMjcBBEY9l3wTdE7Z3l39NjF6U+L
SisQ/FpZcaKQi+0BTVGGp8s28fwGeHMd73Ch5bgWXhOcnl+24/faNGKUN+eLAOUWVOv+z+s3eMJC
pX+vkJOamC6bJu++SE7wceKfYJQFU2AXkL+CGh+YTitWGp5wRXCew0tS1ryXM8Un3z1yndZojTeH
f26Mwzf6y4BkC3ci+RiXaa+1WgSqzEKdMByPL7TPWbT6/NAVwXjo1C21p1y4LIEQmaLhJklan6w+
uOFuvc/Mrla60rZkU2igZVzU7M2QF8yGI/Ob7RfXhGJPDad5IRGGgOm2/AmSc+u5bXhsJwACL0sk
tMhAoddTdD3lxxvsrJN/C6e4EyzRnin7HnCk2TC5/9m/WFZ+Hr3XKLw/pmJh0KANbkSFJTbpHE6V
Dq7k5Fbeu3L7rchlJOVY2882kOiwKM0sHmGTTsZSRPCmfNJTYddIkaSRgRAlSF0zs7uAo0+yg/Tx
MeqImACi8/GF+1X8D6c+rRJQUfh6yevamOqWmNRNC8PBTPZ7cKjh1tQV0uwEnTmP0o0vb/16j4DC
xody4/2GLx/eBBi7VVRDgpJBHHj2femLVSyxcLhhckQp3SaqS0XH2pZCtb6Azk/a6bKccla5HrOK
PM20icCShVStPyemez6lPPs0PsPIFpTs2AHzWR+SQDQoxjhbwVPBxxLYraAS0NVwdgobHinjLiHL
GomvRehRbZ7kTmWux7gCMiviZp+qfeZrcTNupQ52UO3zSdTs7Z6GS0O2oS8+Nr2qeC9KnDR0Xv3Y
0HKb5OmUwNQh7o6cxvXuV3crA+MdHr6mvcSQTl4gP6KL1ocloWjVh1hAV1y8sYPtlNpLVTUH8ZVs
RFyEQG+ZXufbZzL6SycbCthOGB9b74tEeqtqrWM2TOHVZc9X5Ap13l+17ffLQ/WDebjEIbgzqFvI
ZOqSCKXyC6K81irM20yTtFqG+IMBwij4VT6uVb41Ugrat9O0CoFl+a8zeQjZcdProvUvZLKszzUo
mJHQO0e/sXr2AoH/csdnXQQvA5teeNo7ins8FC97ZqZL1HkslHVhYFMWpUlnv7RnFqZiGrKZ3LjM
yOaPrQ2IoCnFG6hcQ//1q7jbgdWfET2OEMYkzKxMN0dwkF3OanNh7YvONvrGWQgTlQtADOprJsoo
r/c9JDQuOUiyUolo7z3DBcRYtDjl4nV0e5/H5ktiua/9+0pJJH8C1OcYTbJh7psP3Hz/+Z/QXgU0
jmwPRiK2P9Pmo4Qs4yKseYG6qB4vU+VrKHhFYLaQba38ZHPtKQs0rxV1nNh4FRNRXcOADJwx95Zk
bHt4iBIhLMmVutYiqMZJiVQ6LEk5KFlbCf7vgxUN8C+4cDWTM2ZNHyduFZUGE3sDhIRG0zHr5GmC
Qj7yJ/JPHLeLX+Li69BfEsIb2Q0bQPDz0GDtapsKzqhX+sEhZjhmI56PiorB4qIHbDg3Dk8p95bx
v+udAkuJJa0sOm5G03ZI3Ou+io7X0ESDUMAs6NGfdpt3V4PclJgCiP9Gbo4sy4XgqRwdPEE4m/XE
N5ls/HdgLZ9l0p8gzsMx9QdOHlWdFCZA1TplJM1g1WcjlgC1DAtnKGCFbYLgbXtYt/XAcLJRgOFU
J43ktaCO/dS8Qi0Pfl8PXpRwGi8v4cvjGukobMUpUWe5b2zreFnGLzD5ooJrvZVTE/DI17GO+1Pu
4WgtlDSY5OhUGYc5RGD7L2hf29OMbYEHASToGqFqAHy1PmXc1I5ll5pGTvtBBo4AP1SJo7TMTrX4
37U6mut1YwcUTjpAe5LCZdf5BRLMxKxO9SlvTDbThcqbZ7ZlbJqUlTjUMFuopKFwRufV5QhL0ivN
hqo4RY5aGEDxshG8e1dhKP/AW08oZUGAdX2Mtv3quUO2bnOS4oI+OH9EYBI5UjU4HsPGO/JoiqUG
ALqWjQqPoSqsxV2gP5/NCHYTq57mH+2jXjEWxMktJ9tFTOIpKMHUjd3/os7WCG+Ab0PzqJ8SiavA
h4yoiEWJ5+E5SYaaz9/uzbxL5q00ipyQT7G9Ww5byg4c4bhQrDYWbbKLXBWtM3wNdGNsilabItsv
RADhEV8HyPv2kQStzfyAurx7zUDpOhtjVlbmf6WasAVdwYh3J3EoBQpeOAJnCOGTRPj/p1um0Xft
oY3Ag2Ek83HWbjkjETiQceWE9YT0Lc/svyd/Vpuw6zKUYH5o8LkrkIqbTme7AqXlxEmgQBMc8ZfU
LCbMoNf1mQUfa5RcFGYGmUVQp21aG0pecgBR2h66/mFhb2HmJ0HQMMuHIEdoFFz/IRbdDrJZcNVk
1tgXjMeFTbfaaEqHgQugo/B7oHI0k7iaKoADS00kJldiBDhlEZnSlzdn/PfkAO7VNh8Fj5YznjSI
udeoaIUX+6yAh2wOD1IinubY4oW06SCwi9kElPlTZrU7rPImHcURKm881AjBNmZx28FH15tH0eJ0
OqQh7SPwG80PrZlZCjwLh1Fzrwo6J01R2jqPiU/5EAdRnb3Np/lP9t8Qb1/Kww6mc6PhPUcQ/o/a
NHVcbSWff2DlgE2yTgTfJR4WUck9l5rgCZhJJqfB7Pngo+VHizW5MGSDqOhzD1xJMyEk5sXVEOHx
D+u6Jfus0jYjPrquaYb8EsqvROmoqwd2FSQIzslhfv3Kw94SN0QlL6hV2KgGrJuFP76qjnXcR5UJ
lNwdAKV7YrpX+lfsvab+g9bbxhBmZWXIxg3RTmVr+KassalgAlScDgsLjM7f62NScgBJZkyC22ze
wytcVGsr0z8REeI/JeKu8ROv9b2Fgldbe9jLYGvewoFtixWnIdxJqLIGBECHkQXsjNV7KJnO+LJK
BuP31GXICPSxmP5mNb7lek9xXl0sSMNHVr6WJBAL6PU5CYOX+ETQOO7U4DgQC5rZUZH9Wt2hsEmJ
xjHyWOCwMhfExUA4MycnCoHZa28Y5UtrR5KIYRf3QO2WcgBqfXo9pgy4OtqGp8VPt0cTVRrZqd7t
7taK7ojEImaD+EtwPJjabQ7mrljn0JhLaWsc2lEHyjV7+6cOzJURCDEPhioVxiFgvcoiKbr88H6M
/LE0Sp6IdbOT9ARrGISeW91CgHfBV68heGO2DuSH783X5+nvT4qKGw7jUJRqk4Qgerd6LSd5VLjw
PwFx5+NampwdAsHWdMbgLUxBY32ukh89tdAjPGvrd4LKap2nZoLF+IwicGG7i1XuaeGIHQRy6Z9B
3bkbxL1rjupNhmHCbNSE2S33nrbFVT1HEIixBoM5iorYI8amfPiA2mrL9huKNYR9Td/5XwA50If3
uuatkZ7Z05rQVrMCynbdEUJlvYpsNUDKuGN4ZfWHLz+BLkyze2g9RALq06F6SW4wl8l28zwoJOlY
f2MKuCTZaFXIx9VlUQC5sbN1Fhu9+MQaSg2l63nbqVjfOxSmbKmpDrOWFEomMqKnESGFptNj85h+
8xPSh9l0rEilbWS/erkeVqPYLnSu3DiOxJbDqup9BbB8u+3TUq0abl83ewpdnAsdR3KsENn7i0e6
29mLY+KEhO0OsNDK4qspXFvt2q6J80Jdk9oBcPeScMe7ccL5kPZKLZHvX9rjl/MKJw/3HVWy74gc
VGtJMlSuO3iRVErYw5kjsHRGQeVvUzEeY4Mp4ZSfwnjpZPhj+C6yR7y0f3ZWHTfU7UnuUGhslSBO
8tdivNZQ1OL/chY3h0C+kfJPz2T8af/w98a41kG+eC7F5klxMjuFy3BZNgPMf0QLkmlthhwfJVb7
WK6872aNv6ehgUVbU2OG7BpMpvPLKBqOkuOMl2F9VejbE079A+uQ46gzVU7TeagioUUnjBsHk8+j
YzIEKUWOgLt8erm2f4+mxFUdH3RA6/KZ8lE5kgkw3+ILxNIO1x3jDouoXqYTGn9dhVMhO3S0+rF7
j6MCqNlFhQrUNzAghyq4hkCm7KQk1lLlAHlFl0/S9xOXxsvMNgCl5nQ88lGNfO6ISivas2z73bEA
/AQLKcCxSY407zS700sT+4ckr5A4pFikD9lo7ZFkq3DPIfeYEOn1BHonb9vAJNiYH9LXubqV3z/5
u78/wWkqGZeFy/DYakf3g3KpCoPWBMxk0abEwwkQKKTo50ydoyJaHRgp5RDcSolgrN9h8aTjDnn7
2D0WAbMc8etSk17SkK6yHE1kBdF3eyUvOBcgS+xyIZtDR+o2HA7iWsakSlAhlNwcugLyHHMEqEc1
09knaN+9sGvyStI0DVxaXVThv2Tj7zZyAFZiVy8DA2FQ2V1jfiD8EGOXy0H0mXG+yg+0vZ7MQ4SQ
SBlG++RQQxvwMgk1OW0ZnfLsHgP2zNmnbj6/qNOAo7va8FgzC9LShbrRNw9lxsu7BzxsseH8df3Y
brd4FcI0uhKU+TM8fJVOcXhH52DyQpDaGvqaQQTsgROqXhRdzmT7nJFDiHb8EHbYG4ABB7RVXc2/
/tm+rcO3Zc6Fuhe4MfC0XbAVX+YXl5tzMcr4nQoHXt3kqs/K2cUX2pnulYGlkqH7X1cVV2xnsgKm
63VggQONYh6oaiIXqb/eye2DJOZAcgdnHeeSnnxFuI4hiQVXY5a9n5bj6l0jlFG5a+t5OetLGsp+
d6vJ4AsZCWbc5wGNW/xLXI7NqNekpT4Qw3oxYh969Q1VOiyDScp09JaH8GreaIaObIljxeEnWQaR
RkYp/7qhrIaxolEptUcHg5J94kWxgdOPozBVXNMHNjkWYTgE2rLKJNn8xKbnEaLPctY5FhTE23/C
hQDOs8pNc8ZWqNFhQxo4up/vHfW7HM1sRVwB+uPy2dsrohxfI96Is14TgGNrfwo64D2eQCsSXeoZ
oRx9vD4xAM/DpEfPLtoaFb+O1L4RSY6GrQb2+U719SwCKkVyNcGXm/I+lvX0mQRsJeKiiEe+d5E1
BibxGo9kCtRz2Afk91FrpZpcmbxnbj7J0XBbDHPFHX5zkBXNF7ZX/Atw89kqtxqdjb57IdiiwiIo
XtqKyYuz3CFP1EQmCEBUSIf4e9/cgI5FMcatddLpV5nUbRHRP1Pa3QG1QwLCaxQAIFcOEXg9vXuy
hl+fJpLUut/cNBOnUfFeS52b2pxX5VTqIMaI68l8A5HVIlUgJg0aNxLWfzc0famwpY7aPDI2T9rE
nKfvtkWq+HZKOyOCkwnZ7b6xVIi95CK4fAma/W7nUoiOOpVPNHZZhoQINHlkQrNbGL4N9phlDYyI
awisCb9UNA/EJGauXZRpO1IOi+0QkBz5vfiVAc7LXYcKe4SFt0ZXBi9KMrWEClIH4K47mXHyi/Da
O+vUoLQ1bQkE/+/stecDNRAOhU6iuk+y0G+58fmkYSsBR++I6Zxjvq+N5HniqNor8AvwrcEocVkT
TFwE9NYptKpFZRv6Pw38pxFa+oe1NCLUGjiCmne4IuuTJCNLOJnXLiIJ6fU3AuYWcG12Vg8lSKiW
DLyz3Z7X2bdGBFVMIbw5moiGzs0pOfgSHxuInvXhvrFSuvtS+KKODqZDLdnXeDGBdyM9wDjM05ro
Mh/TWPrk2E/k5RhdNJs8pA2EntXG/aACpZ8iar4nnPHC6TLQBGc191/6rLwOwA0pNdnGKVuVe1Jj
l1VlFbLVgRAhAvynkQU9mr+d9UFE6u9RL7Ag1KWu7+RusE3+Inf1BzQS0JWuQ/ECdCicbPTXPmG7
re5hgk7XcR2XTUbX2ZDdejdXqQdXdMLUHLkwJwOcJ7HQjuSV55RVO239HtIA0awdxBq3rsAdJByW
awgn35lnoCP9u1jGov2tmUK5eQNKII8LAkRm00vEU+ovliQitIQ+LS+JGRqf79buNiGaFgCghFaB
SMj6+/WS8mRwRaPgn1nDa5WgDTJaDHmYgn51Vp8HkW4FihG24KBQTbPbmryst/1D2pqgf0OD86wJ
7webyK6clNDm+zIQABlkXFbnDSdiiw4OnJHo/Nvbg46QuKuxiEVVzlhJgHC9V4o0TCh/Mvt5JJOa
hKYWI33hm4fHz+NGiLYGcnMkNtLi9usqW/mUknZHbFW3siAxVSc2LyAfE9t+I/LVZF6ATecXr6mz
Y5QKs/kVzq6WlpPTds8oFrtQ482H++Oj18Kpk+0iNWjsrvkbReb52FsFfLvwc9iQqXw3D6L1lBAp
KV6FT+61SJqVonBPO3F/49bQ7efx/Uk0k6cY3wGFx1Eld0ghLN8/lGah3NZYLDUmteRg9hbOvFKy
X/7QYejObsfsdfrITlbGj0c648ycF/0MLzHX5V8CkubdCO4rT/vCtEma9ComPCpQpYGh+GFDYtkY
h4s98fDPZJl4ZQylUop+LCcPkvtrQ0zuWTd613BU3sfzhE8c0Q5y3vkuqtXonzBmqqQbtAYHbggx
np5bUyIapAqDJEu2GXXLneIQb1Z59IpOAqB9Mv8t5cvf0lPhDcZww5DVJ6+1y9RNTyfHRs+243BE
ZPhbalZn/x9pHESHhrq4Bc3CvXdIpOKEMEitYLt/8MMXb5lNCtR6cou3r/IdFCiknpNQnQ4or22Y
bz1x9o7IzSaaehF8zAlAclYJKgY2XqMsk4zo5lNji0nKcpWdq0vMKNOfe93tZqeVAZo6oEq4ALis
8thUm38rqKM7Bg2C+pt1fqlEE2cVgRenyVd7dz6N+wHOQhwLlI5chLA2rU2uqxm2lC9sYnSoDU7/
w/JJ161aE1HKpUYSzJVYr3jHDBzECiRiopfVV5eRGUBNeC8bnpXw5G/snfCq/kriDds++OZBOlbG
+40tN6S8ED2alwptcoBwJRalhX9BZ0hM+nWx7MvjrnhMHv61JizBaCBhGeBf8xe+Lvb9CLsDeUFw
0diapt+EKIVGP33zVJUVXKYYZ1gyOJRKo1kGRmcsYsgCVySWI8fnZPe/60GHGTfMa+gFECZc4iv6
tsbyxejVBsX/GU8onsdWVpnWibgZuE9n4C4p8bRubNOGqiZt4jJCot1sFIfbIOZQHlVo9mM0j+QZ
ZphZjiIq1NW3VUwGUQna5GdH/k5tEKOAuVhDFjkFpOR1O+cnLbuD165W//QdbvqEniuhx7r3pXtQ
nFsnZSHHZXKRboB5rHAEWc87LL18EcDGMstHSnpmZlWhbHp9vR8P1WWVqch9U3qjK6tt9Gk5+0a+
lmqERB0c7S5clt/gKynrBVVuN5G2d/vX7L0Kgps7Asrk81LsGE7FHpTNMA5JDR9/O4yCN8I2/svU
iqCknTH2bvT8TQVAcP/BlKxJOVbeknqyTDCNT/ig9nPOa9bElIJXdec9Qc/ezaw0ngDWoDeyQzwU
atFf48psMwXEoScRZtzn5acKtgp5yEcFbTimAWyo20FRfj0qYODswDF65PTQ6KmUIB7JHhiPKf7X
HlPqe9gsqp2hz/x9tJKjnx4cvIG774dxhZYp1jdDSfCvEM22C1g02HPw2SfUHywvyjXy4Qe/Bfrh
/xV9v8SMdcm72BUMsLLr4qO86qkCvjMAGrmHhlInt7twF7fIEQu79ndB99EAs8310oqbA68fQLfe
Zjfi3Kb+pX+HIf+v2yaGi8zh6zvKcoq1Twq74bawRW56xhWCObhMgpOc32cGkVxxXnaVo0/MBaTG
lojHA0ux6j8QkI2ORDj2n/yVRL2IdJUh/kxdIZIYr1/RGjHP+F560Q+nXTcoAHFGmgokvNK+T1Hs
83VHbxwrr6OpCppFAbr+0f3Q/FT6YokhZSEpzEe3Ww9eSrNfTfs9+jt4CAAZBipwLIg2Sqve1pAr
cQBlE5Koz5PrwYtCdMOZ99vZVUAA93cD1uuEvUUeB+Hu4vLDEbZcGqTHxWDzA8Q3Qny101xFaiyp
rTrdcEP2GRoA7lD/aDp29hqJGGfjrubsrOrUFGEEYa1Mn9uN4Tw51MCFtvRuO8V/0Oq7ytZ3rnYx
GRafsqF0+o8eIX/2kdqsDCiWvuLWMrzIpSwwfX2W3TEG+Y9p3NYrZ+XBYxgUarK1dM2wx2u6vuwE
ygQ7f+DHHPmKNnmBgr8lLEEd4EPx/RQu/OgW1kYvFEIdWipG8/fq9z0sRqMU6vATyClb2RcS5icm
fMddRK3+/oSYGRWOXmXu5/XNbPPhN4HuiN8EymlxVYjRcMQMNe6YI8TzxXc4NX4PuAh+2Da+pWyp
9qFAXLFmywIQKJbbwteCNsRlVsgk0aIjmZ83iKbREUQL2Cm6InyDY0FpzPN25TPqz2n12BtgEyQ3
qULnvv64q3gI+QFB30iQ8PkEDgqPkSz3Skwc5BCSPnm0dZNY9//M3t26TTpZW3WnvbekesJqmVWT
oWBt4xjhykVBWT7nzEYdHhmr1Ekl8qO9Jwp3xgP2IHoaePDf/qwrrgfrNap0wHT0tB/KbhJWSlW/
jBu0nUpNBiQz9QFiQ0ySNeFsVCjEf0TRyidmWtvqqSMs9ikI/bwgolLYJ09mj6jdhgGnLxcYZ5a+
5kwCsjK+nb6SF8CXtpTZiGDfXaEH1MQz33hXDGq2koiUlMASFbnSL36sfBLeNBuYak9MXPir0sg1
SKjGUATQuVnxTMXujuWYnWnUTTnMFB+w9Q3kKR3T7moGVVgAlZ5NRHj6SCfChi5ml1MlkM6j+ljv
dnDq5yCBo5PBG0K/YVdo7JnUK2Ppa0MmHeeXudTBboRICSkrmyJr5LZN5yJHtWE46JmhAq928jOt
eAunTu8WuNqmlc1krydOJyEfYs7+ixDchOjZwR3sNecfex1OOdSMBjnZVUYIhJUOB+eN/3/4I9ZM
YBklS939cP5SA7fV7+oaEBW7VssJ82CzzjJJK2FNerek2kRjKdCnI0+GiJdCYlbECWSImNUL1Dee
dAcIy7brNkPoSJAbECTCoqJU5hjSuvLbrd3x4R80OPnZpkFlK7y1tu4Vs0Z5sPfpf4PblO93lNtj
6ZCQ1Edi0vZevHKKoyt4gqEfidVNYfUuCRzotiKwiYAONeFi8wEY2eNualJ57GPuu/RbnuQfFcu8
HbePwRE6KjgprfEP4RzlV3O1LLiS0AsFHhre3AkSzOaq7uRwQtuqtaqXsH6pOIEJahnXu7w4W1+N
Yfoo3LQ1EWvFg9RuviCT0MQOlXGOOsoSJh9pIqCurFDM6SfPmqpwC17/O7BCD/Uz/Vsq2V4VNXnH
HE2q+2pmYWQd/2Zc6aZVyrA7rPTeQwywQURjlFolqrUtcnzW4dzXixm5CZwkGQCZ3ofXsuJBWDVp
bvIlfgdWsQaVetSie/1eYzULOY+Zz2PLaOGc6xVOgKe1JE9MlTRrHhICtBZBbNfrVoCy9pZnhtSx
e5BhiWJZ5HZ6stxi1dyyng/3R9I6dCQ9uYzP9vAVcE+H+I3KaGeLx06vdutfYcj6A+/h/BUCfJQs
4/tHILLamyt8M68SmulNaxbdBgxtWyNUjhlupn3pnr9PK8HIFyvsTjHK/X3wys5VDgt1jqfsdC6U
lKugV2xsw3T9DBh8AJsH8bgQ02NWctyCCnUYnC1RoQeABcaaaWRLGRUwcuwkvXLq1YVkQhKZYm81
FNm6McUKEIL67p95e4FTsy1XprBL8MWamqEDOJ6hrdRmh87pQkJRW0ln2XCziFlM0/UbcRWUwnJt
la64sc8lDwLvWXNfhsNaZhPdRL16GR8cCWReHGy/+JaWJzB8PwO7ZNBmYZBIDbB/HNXNRxgDEdPO
jiFNy7sS7ebj8XZbZ+Y1fd7QLScdCyxEGGnaXY2z+lnYwvCRqe0a6fJO9WcdKNPG056MryQ3A7GQ
tP3wQ78KwRi9oKC/3hmmJjsnuBnRQGNeek8n9Qq5SZmXt9J5rEyhu50/Nl/M1w8Sr3BjU+uwP94F
jeJTPRBHZPyq73m/G+fPnFpj9y4CqmbSy+YDg/35IX63gj6ge/nsdoScrtRWYJBvqqodhPh5nwpg
MNAEWe0SYD5QuSNNRjkUGNFq07Eo/Ni4LNKCmeVVD4qECJegMrXq4t1+eK9D4tLgYBgWDaUGqbEL
ccwrYUnEmGB9ACJrZQLgzQQ0IZW+uRSi/hwderB4KOOQyYe00kgnKxvIWv+KvA1eVWG5+rG31wrj
KRYL6AK9sTN6LohB+HYy6vnhPn6OervbsJ0zsxmobIjS51TyaeKwVQTCFaCe4FFqdMBbfTJrQEgi
J+vHURvNfej/Vl3clFQ0kbBeFO+OsfvwkelB2PqcQCI2moZ3pMDwsBu0UhfqTBcpiYUvx6Plkgug
aAX4DXoNnqvCqeZjqWZRqyoC1ZpIV3hlYaMW+XixmgfPKNzY4F1bY5I4YX9nHUE6yYms0eMJF98T
TeywQy3bJCtUlzFIwnPlN2Qw8k2Ko7A1ZKN5lLMQmytYFopZf53vJXjy6gc/xDnqoVtdk4LH3rhY
NTZD1WS3K8kh5sA0dqbLm3PgkU6/Fb/wHxSf8OepvtNjumqJtqc6NWs3g3NRnnwxd54ubdbJYCio
2EPkqpC5JEjQG3HqkncqNCEc6Tr0htBDTL4nnTZSK65fGv20e7F395rA58qHbLkSVrYfgKACKRCy
9ytC4MgKGB6NMfoC2N/8Fn9EZqGoet+v5pSlMeU3tpC2fjxFFG8Cx8b8dW3g85YfyeaBK+fxUSR1
0LvuorWmArhdy+IN1/Cg0RdSJxABG8CSRghv1gghUaX1zia+dq1Wm/a3qzC/1h5hwT5q06wcY0VH
vV65syPZ8VhP25Tk9vlBhjTzjyYRILzaWCu8Iw/ZUg2gZJKjQu27aHgU4pJVXWs1bhGKTd4W+cqS
Psd0zdFYRAFGrFlLHR1b9zjIV/rkCgoTrqNcJTlpiewPC4iMu6D45qaLK4vAAzewMjZ1GPmMhGF+
qx6NMnZxcEE8Lw1D3SR1hVKcAOFf/ovBO2l3ofHn7RPGf4+EoavBjrHExY3nBo6OQCI//G7rwWCi
RijjokJ6NRAIqz3BpzHZAS1KJo11ZlvNr5WrMq+pJA+VvM1S+QWmYbntVDNFMBomoSXKdJS2dEfq
+/ONcoDQnfTmukVFMb6Sshtye+bm1pDlB8UNurcVeJk9cRVjtDMKEH/u8ci1E76JiU2cERHzjd1O
a21gc3z7dxFalLyxvts95ixNe9EkLSz12OFv/T8Bewbk2Z4Y4oZZrnzWfOAVSr2FVYSFZ1p6Is7A
V69nrZ4kguSGd/Bt1JEj5pieKBoM3WMX+B4JBVtU+sgOSycSNisR7aa4wkfuQiCDtuvY40lqBT03
3t7gN6Yp31nYOoiL4yUAwg6ca1//Q7/LUzveJ/miXeXzBQ3m09MFxTqJqU3ayGFR6YM7YRrZDmUJ
SxQSBMVsashkD/clm+bFthXYNHdwGOrSKD395IulVoPW7rInK/3ttEJ3p7byRaj9geCtB7R0xghR
IWPIdX5+C8D5wp/9IxBAaO/XGao8raeg4nxvfo1tCHXTM+pBAxU4dLK2M6n+VyYS0bqE3QuRWTi3
OQEv4WqEpzY3h0wJO8w4Hsvj1D3xMJMPQSdOlUP//GNpFr7amZm155QV30xMyT8fbE4emswtCqv/
AyMmDL182nPa5G1GgoVpMBOB+MXfMvXZmVgt/6Ya6b36E+fQhkJ3xJQ/AJgplqxjU6d7srS2A39Q
YrR6JqbVH1CDs+VSTi860RacpPjoDRzUU1Nt6K/HyGOEUrwsQhPxWrbU+fBVs3Q3LQYslkvBdo3z
qNDKi9uY/IHuIeR1B2dDqnYnlloDGJwyhHUqqKeNFy2sjR8MRL27OnpMvx0saVyJCddYklOEx8L5
m0EucPCIEitykqaZ2wTNcrUZXkXNMJVQNa6TYeuhN6FT4rDSzXmAJWNp4TP6LQsjMO6g0SFhVVxj
ZMQrN6MSAQxuRva2ZtUUWHcdvkxUccD/15bAqRc0mhuQbNQUOtVCAYX2ZzS14pXauAxOGZoaDbTW
Rjcz5utw230UyBIr6TmV8MAM/GeHBHfFfBkJH7laQ0E0PI9Y+bqFmnlH8tYRz0Yc5r66+w2eurSr
E1YpucDEHTIr6TgrVWNWagbkWcpWkRytT7B6XpZS0Bs+6YXbYAmk6VadtOZBG1qMoAP9eUeIsBJi
WP11bnAM7VRDllWtadVPqohoVkgDP95r4N3ha8ykkzvDmzwrJdFEGC9iFI6w1AplXBSfMphDy9YC
pF+Evf/BYZxthA+Xng7USq0os7twF4AO+c7d6BUsFrK+HFp24nGyZF2kXURRFD/XFPTq4OlW32GO
izqNkkx7e2iP0n21V6xuJmCVlk2WbcOLg/r937u/P1wVvXUWgGvckWWzmGL0rN4HppibGrL/VRQ0
tsM03pn3+ni1sP5JiMswwBBDwkNRX/+ccttmuPx1R3LYWFhefPkV7enyiOXDUYIeCMKMnhZgplfE
jUPGa2MJpQ7wWLMrIWTUZ6Wbbcdo4PvUf2eCRKfuN/K7LMCRWHWt/f3Mq+h2qEcJlO9I3e5A3bcF
hZIKh2qgpArqrnQNV1Sh2VuzQq92TvY5rw/+7VDhjFRKLR9q1uwAye9Z5uA+G9Rqh29HJuJrRjhV
K+lSbUDaH2WttzqBWvQzM+cpGEgWsqyTP0C3ZcRC9q9nIK1uF9rU6DM7ku1uf4i23sFqXRU60UQC
5miuMfiCERrXUudIGauTkQJy8r5/1Oh91T9PJN6i/ejWe2nFN6eL1UUvhgjtThhs/OqJAcv5ikWe
mdfziX3p9D/iRERFlMoU7HSpW51uxzZdg1A1zmAq3QL+Q6p/ntX4EnBmwtN17A8g4GoQGSOx3jm4
3sTHtqdK1D4yo16jZ1Yn9zI1xSyuJz7E7ZfitiwUjFOq9G7juGm9TcvqyXkpA+MnJF9KJOjgk6zf
WjQllCt47/f+txP5g5PCCunrG8wTn1bA1OUQ1u3J0mtd+9P90MMjqNemzqnJ/OEaTDi8ci1tPfWF
XTdGo1YGi1LK+7uizmnsQhzeKyVg2rATd0YZnrXuEGkm78wnn2Uhs5JmAL6QLA2os7FFG673QmRM
Ufn7GRqC8k/qLfa/J6+BTje4Pd70pOumktX+p2PAK+8IN/Xyo+Tx1GHfVsPxCDYdkxcoGOW4ykhv
WNDoQ28nLFTUV0D8ViITGRBak/JznkjiKa7Xu1y1eNJRVKzRqZDfgfhk4p5VM84EhoR1zCuZQ5gv
4JFWUF3mj0DLVU6eDduEFFP4s94qeAfqyIv6BWttQfMxb4L05LQJDHYYPU8KB+LbW04HY++zObsD
9T7GTFVIrev8HYybsrbGtZCo+H+wlb6XpY9aE56S71lNOmluqXPe8kNMwzrhWePhqIXIrfd++yRP
kyjg2pd7Jk0tplazSDl9wnnA9z7XicLAil7xCWmmGSdnp4RepmJfPRBeTUusB3YlbODiTCv8Zbhz
rZcVwhgjIGYuvcKdFFd/ikpkbAD7xV7MEtAUpsr0mYqC1V/zkfTUA1KHIUzAEWJAWI0SYpZtvpf0
XljtLR9230Z5OrPPMK3IZxq1n5G3rid021lMXxs5cb5VTyqmH7qSF67ScHp5GWLfbxGJjqVog5lC
ciujd2jzskBwXVgeisTGvg/y0OSxHrZ49mMASPaVRpvfqrIbdcfIy0Xr8gFFl0oZPUu+JTPTT8fC
/hvx8PsSnAfKWV0vG4HGJE2R11qsYnQhFNl4r/9sw2YAG4JK7Z4RWgS8fp7dFNdSgWqKvOIFDhvG
c12z3bIj+6keoS6GLJg9+5fepsjfFR26ShA9lt6pCWwXCblQ9EiUQzq9BsyH+9f9HhGmXO4gnzuf
XOtsXk/XPbX1k96Lm2aYASy9Er2KCH1Uz0fg9xpFyOwgbONOC0+/VK9PQmmlAf+SbinR++lpdZf6
2Eep5wF2NnzD5yufdSvvXeyry3Tff9gDUZb0BJOfeyJJ5Xww4HK+Ky7h1cC3XytxufG4fO/Jqkk6
+zqOmQiZzW4uTvJCnIJKHhaLw5poTvSb87DMUcPYkVTgyRXf+ns/qpXsB/ZfEkMOqbWn26osSiOc
QG5D3+RrAOXrU/jddOOdMDSwY1o27Y3fs9g+cxxVh1DoSjgoVPZdFWnJiOFN8P/4TN05/2Svzbf8
jXHNOCvAdPtT0ioKNyZQpl6C8gok7EYMt7h3MmH5gN7oJH7u435Lec9oAfx3vl82rJ39dOVHlOv6
4N8gWw7esRTrjt9rpiSs/np19nMGj8moFV/plTPRplW7Z4pzESzVxCwH/tFCHa1cHHRuvg9vsHed
P9q5GjwARoDywxjaTkQxAGp1A0Lk9i8LVWbpnEZqi5wX8TlMsBI7Tb2ltnykqvjhd/QfktX1X4lW
4iGxkkOPlW/iomDzUsexhB9n9sY2aqCu7aGRozZFvF+KvwQQlBNhqWp/H2yun50WIzOMa6/vgPgv
hce2LLNKB3tcxQhClVKWIRIfjn6N1fh+cOhyyYpbsaOBX+7X0FodEBQViqiIefSnhQGt4as63HnR
wDqqzr3BOPO71LfpMV8ad4RCMpfekJw8ISU5gqAIKsz025iDxJu+1rcIAij2fTm4zwXAccydmG1C
HM/VZ6IODGvC80TioLaMq8LmOU3HIdLgGIlNCOvL6RHYc2cGWMGUNpFp8+9AVKw+Cz79leknMTQh
SpVfuS0oHxaeVcokzyT2/6u235xLVK+A5dSEzULQXYdR1AMBDAMKZCXwuPhod5uuDKGBYa0/j7l/
uQoWvlYLcUgrzNzEEytutcVAFS7OPHExlEtGCbX1k6+U27nbxSAufiePILS/2KY+CcWU2QycSSyj
CsdRlMRxHoQpgudzFkRwPWAA3rxcnChOAeikdtmbiomTI/KR04w8PeVJcBXhf5SWECM8YU2Xahml
NaW0/nDtvuQflyIOPstm6Q4dHz4L/VlcSMctAiuDmyXtffnU/9t5hlpwP7yLm3/rDJOfMheC3lgY
WVYDc4mklTN/4sDKjb7Lj9MqrGTh3+KD5F+x+816YVWaCxp4bD+yIEa2XiEU8SB2oMndPLF0crXJ
lbgxeOdvtcGdrketgyk65GQefoNkRNSbxiqq1cvkuam6g2x7qRO6c8LcmLNxn+gpDsVzpgh/TDDQ
pFFS5mVybk5fB1+BA7OFQtfeaDrKkxyS6PEPjTwBTUDHnG9ozzW1PRhmJrldo598D7rptKGhwnzP
bzGwV9Ms39JQII2RcgXnVDxlZmJwvescsgx6MgiX0Q8pZbid1cPJ+q6rcAo77IMd0eSbf83miOkN
KCpJ6n8cBxycU1GtQXJ8p96y4r8m5zNXEwhd+2+c5zzNybQ1feGDA0GGAwBWeMsRsoVBijaVh0OC
Omzu8/g656XuwwAZzzFgH6089DYSMSEiiJK1j5pOjET+33XLQDawh1AqA3or7xKoVXE4yh6lXKnF
T41uZ0xQ1H3tqQTGqLvQgxa0BzZtSF7so5EIM8id3ykrCHAAJyll8UeLqK2gpJjY0syQerczu6Dl
YAQhDuw9V/LHE/fCjjqUUKaW/H6pE/teil8/U6kjXgVPm8dY0YDxdSPJ/MvYzZwhnFbVosoqu57R
jC1f9TQ1SMC+0M/5HqKXVFV5jWaNjLMcZgHG7Ip+w08wDjFkUoWdpywAMV5kH4XEJfP6YVvXsZJy
Oj6lAL5BGgFgFwZra9gHfe3GLmH/j4Kr3ppdjxTIMSJDKWrhz38+pbueIAoFwH7y1WGyF6f3erKq
yfACSeq1M6oXMLdQJCemloTQu/te/nfUxbBIavKkQugEmZoKD7WN4jhN9/2dF1khEuuw6Eu3zSoB
raRy1FCfJyrw4W5vhBzjRPL+ML9ynbVRYI63QkClR20Ge48y9S6zhGzWvjYl3U3cTdaXMU22aSHL
L2AvBbAD2291bd9p577LGc8OHddX59BGhuIwBjG5PD6eA9aNi+YWIVDU5XFUwqyfzXQDuRBflkeQ
Axjv0P+7tk/MfifkJGMZPBtvAHte9iCb7uaC57T1HJsj5qzMRFKUmfHnCWC1+nEtAXyOJ5zyfINy
AW3YRa+nC2TFPYaFaaleh3h0aSVq9fqiyDg+BWObERYGH3Geb3cr2N/ib2BSwptWnl5+BorWddDz
UW+bLJ2/SzDw52hhkwYHQdCHPZ/eIDPrLY3s2kKluucjB1CqIcsGgc90G07lDDhOev2SwSQgS5TH
lphumAnnYwJcjvyu9wgnOfugeakilaQGQ1C9RAAJuXl67lUj8q94vArhj1lvQffgauGaAvPYgUHi
rMPA0nD1XuGwT1i51W0WuMVJqaTvzU9SWYDdJAlunclkI1rZRwP9G3GJzNeWHbvnHgajAkTihTe8
RKXbd6nA6QC5qGT9QTYJNbHv3HcB32CMDpe9AhOafpz7GKYUVYRbs6LtW+38eLqd1hlwkit/2RDa
tf6GnE8aCZW7nhbpM2oDwQISNbc3/CN+v5Otm1/oOSlNUdh6bTQ4JI3FzCFwW0nNcqK8Kim16XAN
XqNMkgm/ERduwi6Gp0Ic/NuO459JIvHAw/oYfeG6XcItNjCKh5Cmy289exvJz/56cC0vVMwrt/BP
oRvNc/8BK/CLfOzxZOUpHT70XqkuOWgdAGMxoWDa13/1CNP0aJb7xAKb/fFZdOrzoZz1MXrFrrJT
kIKVGe+dDR3D+2/cY6sPvOppriSFFVon4ehtmwL2EG5R98ra5Jhk8x1nvqI4fiL0DblBEden6xIt
1WBBPnN7a9rZj0UJVXP9YMGm76/i5squ70s/6HL8EHUFRRwR9oBd3gZrtFCxabT0yjrAFyXLWN4o
6qJ/xmlQJLopMsXt+obOvA3lGHdFwig4FZyftuAyigdpztGnzRo0nE6WFXHE05fjxLNxG6/PGr12
iwmahg+VOxftBqur8lzktZW2u/08wwQp1p1b1ZNo1ElJ+KcCg20YgnXI2w1vGvsdiCkuVJOoYB0L
JlG3MVaPrW7ipbVblXqa646N/L9mH5x07anhbdBdaIc3r1NYD5QmAiKMcL5kow9jlK/vsnM5ynVf
VENt7O+bKNqDH9xDETtKbgMUvzf3dd6+GPDyiL+9LIL63Iz6enXuSFTDsNBLR+9sDOzA1GNfo43Z
7tERqG8EPj5MDKIb+7Q5iHzV63VmJJ8bzWz/Tvl+9aLtbkXH01e6F0XcQDML+xKM0pwFboTmT5Fg
8/JOc4/mdMbWneNmOpNwXu8MEs/6hknPKLY3+u1Ujc/obIsrMNxRA8V1fwG4f0HJgVu4eEuzEIAZ
LpCycZd3n/0yn8Vltdt9TfyICZuwt64LB+Rmfor0l05mt/y8z+vQc5K+oE/P1btkSOPJEffK3SD/
ugtgXdF+40ZWvtYIZOZsEA2UVAaFCa/i3GaFWJsNTReW8oqzhPlLPgEbkgAWuZ3Pow4gYIwxFeOq
WU44RXFFvQhE6EzA9qUbk5liRgUqam3GyIHUgR5fs/8rCK5j3putsgVHSdDsqkY7MAabT01VEw2u
phlT5GXvHYMRAqYqJBhxRec8WbeHB7FtdPCiNupoVOWAE9Mu8xdR0zTHP8YaW0uxDxJshui4VTiR
I/0pf2lt3j2T/vm+CnVosTOCCG+N9rzdLZL61NIgdD7VnxmqieQcHgm9iPP+Xb38Q7/XUstmM2Mf
S7cP4m1u+JfbZwluhPFS+q/ctbPUb2azNImwapCOvxUHn1bhVQ7Um4E/AeB5ZsIwwjNRDuRzmhbY
BE7Pf+Z3yFNd35o4F/rO2jIFuej8UicalrNk916qwAecxgxtkxTIuMq0ozOPa3Lkz9RXwqNoqNb/
UeTYzxNxdbiuNxdPSRHuJnGOwv98GtEfSueBcW+K/lmpnFyFvuuwjnp/8Iiy0akp+cV3zyzKpDAn
+mkVn0si9OX3VU7bVbvzLgttOtHyDeBFGXyL9rKvJGuq6WGD14reSUOwPpQKj5GM8irQkrkshbqs
j0KdeALy/NlyjZZkGvrLm6fZpdXnCJOVpfpP4Ua4IOnKYLj4JOwkeayyrKBCdjwGUzt+FuCIy9eY
TyM9diIoUki4rz52K6LDp7JXXLvTuBb9b/hnF02YBOs69jnyY5dP9siko9WNBHF/GoJZqm0+7H/j
KtW1mh4IbvjoJCM3AdLmxQUtEzE0Td4yY+JPDHvGrF+oia/a7BZJ1qhpaDLX6Tsgis+Rgbp6ptBv
iU4ELFuOM0/BdbncgZUevEwugZR6OT3wQ3WHb4Ggen1ED997wx+Ny3VLXCA//kFed6x4CsnEPR7C
XovdyjyRLCFenh/mLbqInPliH+nLoZ+bzV5cmigCtZt5AvfZElmr4Vdxo/F1n5e8PC5vBfSVNony
lFy6KYWN/QwN6fwQPXHqMPpRKmAkBj2FBM0Ziu0W3ALs24pZqfPKqkzgS9FZBEkM9gez8DJwV9Hb
pMA+D2dHLLGli1VioFHGdbQTnrBkRE7wtN0O7M5G5Zz1Qy4wmDrrAEWsHq+Io7iKMkBET+q9nxSw
AdGXPizDxf8B93TLEE/BpuOgykiFCWXU0P1dD2p3Toa5An4ejBOc0WsHhayKJEPLx7GyF62F/l2d
CnX3qBe7XGeUCsUudRQ+qqGG4fnMN2YOVrHYXp9LgK0Wz98WL+4D33JFT88zcDXy3M8Zo+ZkO4MG
LoGBDPqCSq5q4vN+wvmThhHSizvShcyoz9wpT80gCnqsYftHVraklkY4eff1UFglg0fX+kCuuY59
+adOFofqEhiQeBZW7kxtDYmPCjAcfkOPv9P4X9lJS6zwIJ0JZCEm5Y3fjLmFOTXv04LhAAUCQpvO
e5vwkHGrWu+xr0rG+ZjDhL/XN39Xp8X4CVWS96/mMIGHdfRVte0EGbmk8qqJ1/z/96akN31ptFe7
2isI40rLBCmk3Wh8O3wrDVr5ZhqkEF7l61GBw75zbTMtnqk9WLqZP4qSMxB9IAWw2dpHYpV9Jgc+
WZ3nhw+pQ1ofsXckIv7qc+Biiuk9MIwtIzULEmxLboqlMCpKIfJJeArIfLwtu+KNgaqZ1B8GJ1SC
yu+VDeb7p61x5a2WtROU4/aTrDoZPxkfOtUsuOIVouVL/WoEM6FE1zox/F4+kmJkK1caTxqfKwXi
x0cJFOuwkb96AI+tuS4KxMn8zrxkldxWxYRcKHUOKLzMgPQsxsUvLZkeM5NHCUX3zP+93/xhXmK5
RpG45UhcGjf3sj4/0cbPRWSsEC3NDDpy9qN4dCNN7FiZU8gLl2CdzMRxFQ3yJ7e/jPLzPHvlJpK7
O9sKBub6SYSetHTgR8ub0MoY2mX35D/eJSI5FZMz8+mrjYeho1l53MDqJcsIIfXyxcrIQ3pVevKB
HafkHanVTsB+mvWS2oumP9CUy0n4hR7hpIAKOjyUZmwjDcB7/PLeWwq4I6M+oOFANh3V5zr/Jv4T
GElN3EP8U+5NIOhVjtC+lI1D5vJCe+ZPU+bwUeAC6oWa2b0QsP2TPOqO/5UmmyKOFKItHy+toKOk
BT3MwwE2uoxKH7pwI9RWmiY/IOe/0GSAeqbAtJyQCceqWzDTRCsJY+Fml8F6ItSfzMMFIyfXugwA
Vw5+f9J41JsrBqgBFsoSQxB6dPJBqwYWt3ha4dJukZCZ0D7NJR6VCIMMma5jnBlfXF7pppgxyapo
gZX4dRFsFPdeS+MuxIX39yNrD+y+ST6j9xJ1AtBcMrMT/9sNyKVxKhobUFYM9mZQqLMa1Td41lvX
LHSZogSW1CgvCwnAFCFgnLglB52xxzJKjt1YgVt0dCM0gqPOdtE/ePFvLbrQsmZlJED0Vnpq9Q0C
+pncxZU6/LQRe6szV7kFJkv6UKRxEpQST5XMzzTffc7MqNnIfNlnylGP3J7AaAM8IhDMo0zEmYPz
XAoAlwlrVkigA7lFrFs1dLAWdw4a1+MqqHPGNr9B8HQckgC8nTmcilW8fmj6p/eBj9KpvORxJXP1
3enTWpG7W4rpwjPGdjBg85qmgEF/UyTDWaq3paAaCQiUc92GwUf0qoHeMXewiDaBHWGmjWt2isDp
DeXZ63+8Py/NetXSDAZnpZjWF0UpAcJDg39HLZjSUbhmkVO6U+KiydSUEJomwoqbsIWD0KZMNAJs
2aHr8wmSGqdkXdt2VHHOnPmi0BE624Ba7n1xQK/cKZsbK/hS/ah/Ww7qLnK+AnoXFjB+4T0GSEp+
WSHdu4ULelHKKm4AaZmPc67zRyLL+DsBFMVOnHikRmv6+iRQBnqIl03XwYEtNQydC/y3JecEv4Og
C+nGa8zitb1au3JI0VoeMLoZ/C5yn/kbbUl8QWKYbbkZaJZ6PnhwmTmRT+hEuCeSvGMdbn2KhlwE
iqitIMsPl1Tz9w61+X1Lfgsp/gP1wzX6k3yXgooIiPMYDydPcZN6iG1zcYE3JzFBNVaMqA7tnXsr
cekGKcWo6CIUAFFIeWVCauDmhHK9yhBsdqR86hiWVO78AHTuBkH2Pg42GquoMf2+ASQuvr/dhawb
Ohro1eOveJazVSGbEduCWAjER22oZaSBblRcyDCQZenwz1C6SMZq0XGnjpZc5/ebcqf8Zhr5GcMT
r5A50OrRa2XXCQczDjAkbA/SiIjCm6vFS9/R/Ft9jZOFecTWJLokTPf658Ezm0vJzANzj4HEoQpc
8OxfTTNy0t3PV/Leud+ilLRRQY8hJs2ovjDlx2B/noQlw7FzDb9f2u7RxWWeHSrzSEdnwb3GFAZC
0gol3l4Sppi/wEMqgtaeR/Hti0wl6/Yg/VIKGvMAoce8Fexx9i1tw2JVtYXkpTCyErwVqOFbQH6t
xn9mNP/wQfLG7X/DzCNxE28lTrzdk/PyP/Cap7NE8S40+s4HQzVCXSUHnv8JzUTjbftFlPJ9rAwB
HZ/5hcgQVg08Injw5ZGXiKCnBi+adReBlFoINaj7aLhxnb7O8YsAEauwZoH0r+ywdwCUOrbzYL5R
/2GAYvZ6sxPeIJ0L3zQ4R0t9WVM+Rpihb0FgsYM8kKobhiS5XL4oadJfFnYnj/8ZiVQP/gBRubF5
BgLFLVBmb7b68IwlC0KdxIw4oROFQrxI9gQrvhTNI8/UqZezUACb8biAZEUDR8h75uFLnscW21v4
GX3jfs9RSeNyzU5Ed1XU8XETMueXmy22u74yNCYvBAPZqzqv0t+KIkyxGPFsNcJirWh2+vn+UMGn
7bkZMZdrZ/sIjhL2/OhPaOi0OoTfWBMOMX55KJZbtpI9pMxBWGCel/Ts/kVz8iwDuTPI4Xc9R6j5
2DyKwVZQIsXtxSdy8vYCXwah0iq8TgQS672IYhUI+A+JAWtJJsy1KvtIH/omlZ6AVLW7pnYx5xSk
av0Bm3or0uwqG141H85AhRGInYHDq7a5BIuvo0FuAUkrIBlgafztpC21rucm/NPpmQq/S7EkuY1V
R12N0j6jaoE4lhOnI3EvRLk4eltReJFP5C19jCCw81/WvEOWzdyc6iruos/u/v92ftRBmKZtSxHk
L53Pr/7U8rbIMEVyt5UyvYsQ6nD0t4cPuMofO1e5gXWLd4kG7+XyKqt61NhtrWvA97wd880AVxxS
ad8B4qh4tkfYIo50FUg3oRA/pZoySmOo5OtrqsaviVkcspohRY1YImkG/nOVzHFeHC1DrKrs9OS1
0ihJ1B3WRDWuw4r85sMSFuiAsFEtLsclljoiKXYECBQMfnNkzU75JFuvuKvxoaF/hec+C5kXFd4+
62ZsQ9pPtQ6AfOt/dtFrD5QItxjN1cAoa8EyT1peSruke9UcdB4tAxiK481+AOttgsoh7slKamli
+lNMNmDLSA+7HH2TM2IKLAwtUuemiWU/wkXzH3dNcYHDCayLMBXAWr1E/hN/YGCcVlTpyUkV0DSr
YvXg4GzcX0Y3l4NF34YGjrCA2LlZWvC3NOJ+qZ0hBHN0uavGXYHH1JJxlhe4V02RCHsF8oNYkGIX
DflLAiIEaloH/Q4UJQy0UqDuegAo9a/bVKTD79kEnBxChwGjMTNZG6UZ2eg0z3IB7NrH8u3BUCHY
t/YE6A9iPCps0ghQcKDc/ZkHOwsyeCP/Tr/ZaapbNa5jMzJ9eve9t0ZJX8INfvyGtL6K6BT7f7vu
TmXutirtPuEfD9o1RgAFsOxvF9y9qHeHywSiZas35Ec7YaGnm24k1AyEI+XmIV4W4R53WzD8sOWl
T94rtiJOYTOhp2LNpIvVYWLl8XISeV3j+ruqxpLFEByMPowvoo1djmXNGqVZC1jj/eSw3qUr8G6T
xkWR+Qykzo71B5eR8QoBUJwuZW4O/nw5zRrlECEq/I9hhOAEIgPkL+d3780CfMofgaXol9blCpZJ
b/XbUGqiiMzq+C8wr4gAMEJ5qHCI2OC3JxAgCR0apZ9eMGq9j70lHv/mWB4aMLMDYb3HAGRrgwiE
nG7QjOHES1K7EPtp8l7U4lHarWoTMt4+eHOniqSDZ0v/zOZKLDNWVDM5Bd0V6qk8+1IHI2ygmBai
5JnhMGyoyRgZHPBY6Rb/U23Fd6TKIMW+QQmTjLDXg4i60EydqcVtoUXTtTBoZumR5JDWMsSCkrni
dooDLuPQM3sGlas7pjE8mw2XICkPabBd1FGJOR4Bfm7jJ3R2Km+oI92VvhJ3/F7BnsWLRBYAuJ2y
Mpo2+2mMCN073yOTnKa6kjfvXeI0Yj/azwbnJ3HNdKaH9aeZ5DZjA7euvT+h5YE/+tT9P0tDyCux
LyoyOvbyi0TIs+fSwZJJU3WNtZkYOmD4T0NCfsUeOaT51rcBRsHVMxYE0hOX2Tu9w4RMwnsee/1u
7cQXBhDfh0W2G3HAzDuxjFbtVbcWIGbC3JKJGZ1NizgpdvwTGqLQt8rNYVsZbHb4nvRQa78UFjRG
7OXAHmHQAVxIXTVC0b8QReTwtBBQti/7FUEQU3cGeJoJKAuzpDf/lRDr2CKldsfrJ884AevgiWNI
KUXIoOCR/WCIaLP7Uc336fkpkTxNRd4OkprvnFVgI0tSGMnKRQKqgFekizLXTzrbktlhjPIScNcG
RwYrw9GlbXdJBFgzFEdh4N+EKZFnXKFH/Zu2uJxPoRGDRCRmmXRC4ghNwxOdlKbZ8EuV5r37aEbi
mcbreAhVWH9pmxypL8lrhmU/pHd1qTWUMHT474KDNTul+n4y1FMdYbly4WcLVzu790ypGB2qSKFu
FwxNhJICXpCtSMvSBiyoS2fkev9e4x4FT/auJHlLyK/0gABniCD/syN8ddlb5rB2fl5h3OTBhTDU
/FDdc10q2foDz8BYC6vqHwRvKlE2vO8T974IVmmCuEa9HbtDy9jV0R/il5og+F5BrciRMlfpmEEA
wAzPFk0OZT4J13q1D/soTFzKliSluHartCq9imGI0133ng8tBbjR/egbZOdNbtbtVjyvu+1VW3U+
4dWNq3iqQZRFpsZzuQxRQ6WqndGfZjqbndVGKjJV7R31hU2Y3zVTYdiVaZ9Hgvbc1auhgtBqYZEs
RHs30vDO2NBC01ufZCHtbgVl2P5ie5aKFwHO9pg49RC0FDc8H//08ksN7h4+rza8pAryJyBpxVDq
/cEdBI3VAIa7gduteSr3RWrOQchuJh9zxoHXt+kghEeyb9+rhB5Zan0Qw3OCcPLKfva2+MghL4P8
EMx0Mgte/ho+Ujov7YHIOREOhQCS2s2B/cgs3tQA7oDvjcVghbbwBLrpT6YrOmYMWJ3ZAh1oAHcp
Te0uE8yKgJinyevBBWJBna5e6YNdsC8ke88SEqPclMVZk7iJp/EzEP2p/qtpTOLXgQIG74ZA/08e
rl/N8KXINJyRFZ0fgsdi/ew9S1A6Ve9ATG5kKtaukFNifh+kHd0ZUuPCadq7B70WdMCQcmPZpTIH
bP0s+NZ5boO8B7vPD+YRaHXMaw2yo3oZxHAgRpkdHOFsJlqLs73U5qUbhwp7F6fNqZDE9Vn1E3L7
tzDT+tQj4rwCFUC4EevNzEu1R9TCI3GIeOyRKtIlFVPUxGS72U5224RJezAhygc+Z3ipTYz0j8Ce
1tikkxYWrySKj7ENYfeFz1xn3/vMBhcviVeQ7xcEsaiQS65WCDNWumoCuyMk2gG1LyXk9KCtSt7E
lj+5bTSU37OoGTwyIWJ60Due+BKQvuqR/sQACbYsZ4nPWprTiW1k0jxtC+vSOeQ4t0Dbtx5QM96A
/WJZFdaOU9dW3aDT1C8jXZDki8ckn8wzahi6kLYsPnfICd79Z/tCA2HGEDmdqvd+zjHLAk1lMFrG
+LjSbeDnzM2U19xkzTrZHNzsiJzVmiBHIaN8QA2C26HRmXh6ZTj1b2PX6VxDmAMAnSr1QmegiN2I
ByVfd0nnMAWGX/6gvTYIDF5n73CsaC8elwb2DTv9GlKW6IlhlAxmejXqEwqVmyBL2J7zUd5MBY2z
Cltw4LNSlijOJxC+ALHuTFuY65tWKzXwluI7s5Q0iui1791jTYUuhlRHQod1ku/x6xD/F6qLEWCY
eeWsJd6PBO5B3CjVaPGvKGVqnE4ar8YaIhbIRB7HL+N8N2+dNb93s3ayoZASD+Zb3kRBdmu2jYvr
agk11OmNm4vMFpMXB8s08YJU13dd+2Wh2vgcL2lZkZwlskRZzy5IYDANF8iBAhRhwAKpol58QZhH
nAnLSBg87SRliEGtu/2dWIf8n/2mWS290PPznipzJztetjH9e45qP1kNH1DjfBE8ffTlL0P/5mAD
YIUrW2HvCmBDQm+nNaFbMQZ5rJdvn13X4LHcB7STyKVU0pVX6imzNyp8o+LlJ/mASaWrGO+7alAI
pVTwnkm2qTdOwQeJTH9EKBEh7B1bZNAXjQ2NWaIBkEPW/86v+dDOqNIOR4TcYOtpPT2uD7jAyfiN
FAEnH9PxgTPM2qhe9s8I2hTr6W8ZoiygjddSIVpjK1mRXBZh+zvrdo1mXpOcnoy6/mAZbFpykpw+
NNZocVMqL4GU/Yw0TYXZtAmfeDZAPDsLNE+mD/mCKEp/pbiST+esDt3Y76sr9m1Boq2QobiKynsz
DykghEHO9YFi2IncseStHuOtkCkKRp2RaPtuAYjRCURJNO5DybafmcSnS+BvKG5G6/Bxllc5Sn+5
+kPiYEpwvNdVqiv8d04TiCyoF/AV2vQo3oHjw+6JXEBO4BP5k5EIC7B1ObyY+fsP/Dy6GPNFNCnT
9BvwY8amLIJUIXcrqktHLXAPud5yGpKdrQrT1D9GU9D3BGbvG8tThI77KXYfEpsBHMijUp5zOO+1
fLT3LwlG11+PZ5/z8YazDKrOxvH2MVAB2FuWMnkKw35F3Y/wYOdekVMXzpnbN4dxInBwR6WsWj7A
idnObacJKwzu+S5NYRKAmz7pljVrljGPjk6n3S1Aer9Z4/n6vrNIB82SocTm6SZz66PkJFaseMhg
iY056DY53r3R3ewdXX/cZSlqZKU9woZA6SgOoDuds+qhTF1pkGARoIT2fGFA2uIcYvppPB5UKsif
vLXicAp67yvTUZoq2oB1ox3mmE1aaPOdnw7gQl6tzz3YjLk7rolRmpnImsEdA4txxFrpt3z/wHMQ
unsAGdmZjYkbW2yNqzK2YhwswwKNcCvzga1++C/1SDSXeRkeJ8SwlWSQgkDs4Lu/odTpKIZW6EhO
Z1GupYWAn9zMzgXcndgpD7MdiWDiUgAM+NvEBbdjMisR4B2sS/y1Ks0woqnxt1Jh5ZA0bmkhMkJL
lnY28lUI+dfagalnHDw1J6n/aaIddJiJLXeqG+3U0aB/1OdTY3Bbs58KVo2cqA55Ps+F8ln8PTh4
f9s9vMoGmYpTf0NEwUIVeDzFAq6wkU4A39B05OxHEX4Yrxlf2JJkoZc4M6/G+4V7WPRR2MTgaOW7
3KXeLcOB+wc+xF45kqqJuqaB2f3H+Av2UK9/fmxi/VVU9JeR7zlQk1S7Ba+gjQOnOmPy3huR1QVT
J0jNyfdK17uyWOJmLe71FVfHnnnJYnllgf3eOoNaewQYA70meQdorTFeY9/QG1/K8CfGVx1rPVYm
gB1JmN2IHgYqs8Ho8L8snt9f2g21OzCAgSlY6pmKwyK24ZWLFGH5fsz2El4AGAIWgDuL/tDGNjMV
/HHg1vKsz2/2+AAeOkdcgYtIx4CaNFEI3hKo0YhW32VAYw7/95F85h1sPtYnv8Nb4VJ/MCzOxZ0L
6suTMOe6X1fWnzo7VKkFEuEWIXPWR/M/n9Rx5vIvcS9xwrfo3gtZh1t2AsldWpeHx1qbUgmAOW/X
gBajn4Lq2kqiy7RuptH8k81zkwrGaWRFT6RK1x9wrC/DmhIyBM7qOFTM+OOohEP2ysgsE1taG5CB
+1W+lOQsyFBuLRykPZRcFL4U7jkee5iByPbJdzT7di2CfQp8BOgVCxuVvPcw65WTBVBOPDnYN0ja
8tYgVxmo1YWdDWd99fbsJ3m5Gc6WNcAG5aBvlhqr5zYwPSqokmdeFNWekSBmVEeA+cCWJPQ4CmNo
EGQKNR95v9auyKlp0+7q6J5cMGb3MdaEDfm7VkcATcDLPxDaGCLoYSa64O1nyDiOwdbo6JHXKj8A
+qpl8fSdqsKJBZwTjZ9uOjdQp1aDuEzsveQhDjr9Eh6Dmpyu1LuwA20t4hmgy7Igw1QX4u58FHwl
Zd2eBk7DEakVd2+rj1ygeFB7UQgeLhaSA1knBF7SYxVlsC1elzNWepe0z9Nbk63MHPI7+IhKk9IJ
pyH/voXt9HeiGCUdDfvG9n8LImjx6ks42a9C8oKqIDI0Pz4iWEv0uL7CY/cKp9I2EM6YvOxln/Eo
0AtduffeBXi8SQDMUShb8CSgf9a+I/Tht3Ow/fyQzycWsnaXnc/dX7csX3En2uf9OkwqTCmTccMF
HprPVZNz812WJEeLOt0yYd8HBfBZsaOVEvAajIrTKsobfCqzznYzLQAbNi/FWY8RDPSWtbPVNgtB
k3uoLLAHYPaON/XdBdQbfpRsuzYcQsvSnAbT+cMIle6T3uPVNMjAPmDQEEDY4t0XGccwkNPVjvSC
P6K8LwoalfQknPVn0I8P3KQoG8xSXgFjLPU6qYoKjyaGbw/Ridw0Dk2w2PbMRvAtsLdzqwqkshmq
vqO2vM9BPmNkVzVvsspHaR12giNvw4tGhrM65dLFhPIv77F1ycvFG74h31r5L5g+wlX87TaNzc+E
CUcciVgsI5TTXs7MUH6/EPhRym9uQ4IxMDDRAnVdLxsc2WHs6IpmPLKCAvhDW7KRqnXaDBjmYMml
nHhWScNocm2dW6h49XsTrBM3hx6v+ZQ3xkSd0F6uPlQH3LflB1QbvImrTX8S1wsiDUuDsF3/kh4I
ykvD98LHN2gJhCf5i+YUaEy0T1U3DUzJp0iZPiV5+ppE6nNyWOKYjmEFTgsq6U+7bw+capB+6NOv
x4I5UUQASja/par2AVOpVMaxR5msNMl+lmZAYLAmwg245QWYQgHPADIQmjI4dpFNp0bhWVw4l8Wn
6zmrKA9XkZV9lHlfFYdCCJLptDx76spQonIDUgYKgHKH+/UQriu4dA0nI1E/8Ydqo0tHY1gOuf5o
MAbDA/MD001+pGRdNuEsZpkqLftpYmmPoDw0+RD0tnCNr3UidQOCNYIxFxC732UJuBE1IO5iGsuC
BhVxefFPgbX9YIPeryNFg6QWTfNV9V7JuktI2FoKOa00HtE7dmyiSuzAjecu3N+JEDkKCVwKYCOC
XjAbTwXDBct6+CnAgzH6fYTyfUnZOhaxH95OUnFZyyw4k8LNiEL41RSWT3zcrzP4vnSQH3AVwgsD
UyX7CHGc2tIuLgOoF5zjTwZGJ9uiDiLeZkYt9+yZi5JcTZfAtcnWzkzy7Oe1wjw/uQj+U4DaNCdI
oofs6IBEz9+rc3oFtUn/c9CVfbkenjpsmMC9jLaOJKZdSEIYVbh+mS9JNU8/npBbjAOyJmD+y3lx
mUTB3Sj0fNs3sPvfLANkuZC0ZtdyNpih5MasvJGU+JvD52hWxL+lueU0U/lc1pWAR3FLiSaqYasw
v2cjpiTQFMgaB4V91HmHYHnATQGWD8f8447HVo8a3uOSTbz/PYp7SXpqD5HhdKZpbOjmcnZOtbOc
VSf2dGHa5sjijoH8f9h0ugw6wlebrEiGecyKmcPWffpIu2jl05h1WBqz33zn88d5LWMVAS6qXMyT
tQveUE3iQKuxSr/Vl5ZWjy6tfGDgl/xPrkv+bBKUeNS0mkm5QlPtTROOornDEJoX5tKtNgr0xcZg
L+9LykStaXFV4lP0JgymLKe4xBK1Hm+WoHyjEsFSPIyqxDQUTcCWjEzAp7iWwKvhqqx4AR6xXycB
YnxgPAPEPCPfqTCCKn9dyoNYmRMTkRA7srzztyysY+eAkn6QVKP1a/tRbsmcSr+TYyQBcJ9D7GNw
Kb8LRBTGz2yrq3jS1/Adf/TwTzX5DFoah9zfVwvP9ucr1mOj2d/iCVPCKCqB+/91dOdDnpoB2wwc
PcdTalFQ3+xaazkeLNmz6Ald4jHtrhRs1cyAaUjKg7hyw58RxEXQG9IDGNTe6rL1X2FRDEdx5mU+
03kEyJQxuJsTOLWgqM/p8atWBLuul21Fw5WZr8jwITh34pG8cfZoz6N4dcXHAK65w/K8hl1VTU8O
N3mFzro2wlQNKIU/2bNEN2sVlHA7vdmOtqQh950om1nSydV7IGN/+WpWSifAprfhKfy0+/wpBBDs
JFExDwM1idp8ntft3H5HhuDaXwMTHcQNl+STuvlNlD+43HyM2KPUGEAK3kasg5apCjVSkofZClWj
dCQrpqUPazu3/RETJdEy+2zlYxXSQo27knjhWRNQYJiY3fVG/VOkMzg4iUs4TL368PMm83qtt5GQ
EXFF82rPoW63br5mYms6fxn4XWf67IGRd7jR7w2NAsQ0dtr7gi9NHsIrF7ZAFfqDu0TN3Kv0wTFh
945VKNmit4RNQC9fGOgApeN7AqWLpJ8jHUMm5sq1UNlMVITO9KHVR7B4E2CEV20L42MrK0AAuhHq
pJjmNyI7hyhvyqmaX52RTVoEOiUkNJ9S6P5AY5l24LhTDjEKBgr5c42Ivay9CG2gPA7Gi1IxJzpd
2Y3Sy8YOTq/ViMCTszak6cduxGZTLZeuqCIJOqE2LiqCn9A0wLrSD/22gXpQ/5mQGQahRjYsC4G0
QeUPCe3SVmyGma/5eFy2uY41RrbZL0k9TxTvQZUjugM/zMqb+WYCNp6vJJGj8uBjQt5LDGv/7Duv
5OvQa/0nJicZFUwJbdqXRyQE6AcmoyFYO07pmDqgILXxJVnnoPIIVeP1yS4ApL+ZPctreQZK8Ju1
YPGbgyFACUS87E0sBmlBEpHlUAsLbUDREqFLsJHaKhTJbk/ugRXOMpWWe+W6G/bhKZgYTgK2D8iF
bqs1I9oXnA24MkIEQkaIHnZvt/Tq+1rTOVnyIfSctSnCejV53l8sBWS4OTbObCzjY1YN4cI0LUJV
LS3Dn2xPGSG+cnex4FpW67ac03NoLI9o38Mv0BxFBjhagPdGgNEAZrheeoVNQ81AUriXyN4vn8pB
u06sw1OEHTSXSKRG+Ow/ipqaEf8frMJj1V9HposKDcsioke8cZPHLPNaxooRvmMFkipkbBsAg21D
9q+ZQW+XCIBUPaQwfUpXVGgY1vRSmdjOxhUYv1Fq0LtlPzbipwmAMRQ/eg9ttmGGuJRrNf0Y5xmf
8XY8qf5xWJuEuwxcngZ/6hAdbvV8qFazjQby5D8RfNx/OwC165eg/ATmsUXljmMX05sgMLVCUeIt
EyQdoW9djdCLhQvEarRxzzmLsTZHVhQmi1no6lGQCKX1i7eaS5xMcKq9Nx5XGSY/xFZ+ZoZq4MK+
oeVRq748EKOe/JYcFLs07D+t7Xp/+EwLHEDf5Z8rVt3Wdi6VMKthKZyd/kn5yNQ5ozvDU2A/RBuz
BsWoB98DySbda420XpamyGOZaq1QL4UWh+QcXMZY0DTsXaeUTpD4AlCVVQiLwzVjdVX40tgZsig8
Tk9XBq2aJV+8J4DXW+J8uDxfNKBpcRcfsm9lEcmvSdsHRoexqhvDrrwRgp+9FLZ1/3nLD9uVQF0B
NTZtlqPJcAvNVnMDeKOKCmwBWtisShrOa5yrVnWn8zDxr6OgQ3aEfaN1GvDkuCIQlIurgttHlh5R
mmLO93+j8qYakY4nfBPa15SnNNFboHA5R2ImbBguCWgnuie7WBjhwrGl3x6VI8dio+fIcgmYc1iW
AmdzBmOIHRCHQnEyZymWETX3T1TFVRKf9saJbCLghasFzmARjcnY9mzRIOLHzLE6/4U7r2//ndz0
/FiSYGaSv0DMVK/8xzqvc4Ofyq8J6joo5t9u1ctoLqYtN4WlinkVYzdsARAbkjsD5dTsp/ElJg8B
V7V1nrqRg42qqwMPLBpGuFlDPPRmkcCE0I2TGH8Twx3P31MRzllU2pNJZghwg3HAZF4BNU+/OWia
vrwJmn6PpfrxfXJFcJqiUcHJRd29i8lZB/yAkQy+U2d12LdSWWzc33/MESAjyHVLUZ/4+/HMzCCu
DmUW+AJ7Mx5bkGQzc6CLfjJaLv4wjdPAPkwDOauv5AhvtbXoUaCrxmZweQ7K5MryDV9zD0rauIsp
g4Rl+nTuJmN/rPMDpXgL8lOxD2xNEZuoA8X8UCEbNENtFyIerAt1X8F+jFslsPb9S4dwvPysmheU
bo1puAVWA9J0GLK8s2vlOEAQ3tyj6AfCoxeftug5PqFYAHLNVgq/8/Py5db9CxUzd8y0r6LDIjfp
0CXoCO6HedJHoRCEzaBrlaIhGMQwao+iFmiHRn3zY7wlXRCjFxNFJ5sZXnYcSAj66I2v4Ef2gFJO
m7q4JVGYpEw/EAm/hcuNsmddBJRwjcJjvMwI4V2ZeaAOPu1bhVOPQjIL4wqaCut4zDnT4+a0XDWk
+6j/2/NMvIeEpjzsv90YFWOFEVGZ/4HNCq/sMyM8LaiauXe59wmMzcsU0+vL+Tj0Hr6qPn5cdRs3
Law0LDxTcKH6Wo2BytkTeUT8k6IyXzJh6gVFMMJ0J6m/avFbxHsudEugminj9nnhZB+LcENRqDcV
alcRDGXe63pvtWdTUhVoTspQBQLTkwA4sKg+rSHHPbjh4nDGZQg7KifiReATwLmdkwOOjVueKxqA
I2dDZzr5NZ8vWOI5brXtU7/lmq7CNxWePeYmADKTdHGaEKwKdkrVpad1fLBl30nl/8fHNqeiKcVI
HgZjKvsveeWGWygzQIGgbH+uOnXF0cckcvPdHTfMTDJ0qtdRljdQcp6Emkfh1b5eDAJ5gjvdeygX
LJ6Y672qWxhFgzhl+PGpDf9jIrqBNqstJCusErStOTSSxXi/KCJ5iorRdfH+6f6Zq+fhHB+cIdDW
JjG/KStNmSVSZW4DkNTV3fvMqoZIDwpRySXc2ekrV5VsDBi21O0lAVAyF8toEOxWfUhfFYrIQP5v
xTFjt55cCd1oLOd5+M/iOEPgibthhfN987M9VV+isuvZISXDpSeEUSMpHLWBpTdqLIfMUkCKKU5Q
iYCzo8VY1itXyefuv6Eeq0PC8JjzPjNXBSxtdEVpRA83XxGoCMpp1m+pRO3zasGL+x+SHT89AU8D
lOr3DQ+gGQVy7UL4xNDa2hGA3h2m6mjjEJO10bBahRlq4H5MNm+j7mam5hkyr9GOllQYTt5QSYrn
HgnI8RkJZbOrjTPlNEm1k6vHkWbqvKFLyg9Y5ye4K8pRlQhQnY8yPG5zreSwExFtKNS+TukspRSd
SBB1KuugBs6T3YrwQciWvrt3vaa3kjI6emtgw53PqKthnFGkBjB8jFRlTh+LfKGcC2x9Bl+V8vSX
yRFXb30aqZ6srIEFAtvDqt6XpNwQ+19r1zX35G2xGL3T1sQbjORmiI/jvdO0NaLIzZyNDLilNEnL
w2GEDUpsij8Sw1/NBk6J6BsmneFCScG51AGEgITnNyXphOABagrOaMAwt+YK7ymKiDsW6hhn6uto
WAcOzMiS8pD6ISm6KS69qkSgJKIsGFhaACgxmld6X+kfmagqO8yTogsOnehLzyCuXqD+FywoQ9/K
kol+Ypu7MGGeNjgTJA910HaZLgqda3pczjOfBALVSc8COtpiykh3CXYpMSHhTE8KdkrwKnb67LdY
roR/a+HxsJOxthw69yoYY0D+3VU67pdOHkntc1DAPsv6Z9ESZnrqokvcfGoz9eALQiYJav9s863V
Uc5F+Hgzd9eQ0NPdElGZQoN8zkeDpXWhGAtzldm/gvdArvTZw5FbnfDS3szeCDpE9XLErNRs6tPU
yfWhRyULlJqlLFqj2G0VwOrTb4z2H4NfFYOVthLrX0jFSCiI+6aDXr7v0T2F/dRK27KTHUZq6ZWM
VlJ8nV6i1hzPH2ZP/yBbZ7ATACw0nQ6kPD/9ZFsrcCoOndE+xcsNEeV9JTAnRR4f91NgIEx5qXIC
sd9DvRvczLONt1BGVNBaINWYe+32eIue1U/PZgY5ngQram+m/v2I+R2OpawCD2kX2hIc6lLpUgX6
ArlIr6d2CmFNRWmmYExVwqeb8NpoqItuD9+/Xswt6n42lopW3kuVdxX1VHxZNFyXFreinu6Od7e4
dhIAIZOyvmSTAkQRTZClcxw+ZpMdBkdb+MN0jIkqRvaARjWt7+70lSb1bVsgIX/kbXixiSqbIBks
YUQZximxZjIrM6711XcOPLQ3fJ39oumq0vdnjMlqp2pvJ34v7V6HLg+mfPIhcfn+8429pixwqakV
skPZadrLzQzSQHZpxEFQjPyN0TqP5ISdqEytUGD84xuappWrRn+KoXNG1OszcrKbHFZAegDYwthD
OVCpzn8ZiqV85vMTVtCrr2OYDBMPRuICWgTK7IK6rNzoErt3HQ1KU4rN0BjgixlmXP+SP8/jvgmO
WSrowbMnZITkF0Xhyijh3ANn36gYLvU5iKzeV/2G49gsbdXkKIr29ywDox/2IIzUo8ZbG4hj/YwK
kCOPFrAyRkBJV6SE2t2kMFbqeterHu17Lgr8PPmJlvvsP6I8aTnQ3y6Xj3dPEqDsZd1K7wN3x9Ql
b6EsAh6mT8jYK10azOL+XhwBlTOsIR4NXr3DYbYHx6+bvkKKHeMm3XEA/PoJ/pG3jTfMZNLzU0Nf
EnWYCI4kiOncwMkXSI54HVBNuN811zPhJV5xhxv9+GTA6TkiCY6t/xa3BjidtX1KpM/i6B0Q+Epi
pJLWATdUvi/64zct+MNhVi7j18H09Uz2z+hz4Zlu6DX3jON75PxVmbtxTmLsKGoIzopYBDL/7HgQ
Uz4YCV7QoTGf29248MQeckmJ+sDYrJ+BXYoqUPQboTSoWv7EWW0mw33wwxRj9qvaLUXzXMJFsdCe
AJkwiyuJKQGp/ZdDOEizNMKdAKcfrJ6Kb4CUOMdbZ2Kc2LieEv4MxodP08VLelFkQ/fpIvvhswwe
XiWP9WSCpJwyLcoSmtL/iH7gQWNP9XZM6l0FvGYci4VXT4ESiq2zA5x8VzMn1u2de8DoFgvriq8Z
28OIi9Y4c8Uau3FASqcSZvRxEzxu9yFd++/kp/HoMrwxq9xk9Aes/gAEpDCuLaXufVxKDOq7EMbP
of1z5ELam6/2O0BJSNsNtUbmpmGcBgfrjS6nxIttJwI70oXWJvDIjJScsDAQlu2wVpDSoAzR4yY8
7UZJTk7VwbL34S4M7SchImZc/L5xQPMtcZXB7FjAfcf/77c8uf+w+BLHhf/AYglzL1PCkAvpp8Md
/hJErnskc6GUbOhO5HH2lXj1le+TuAMx0qGZdJDT1S1TCHBraiNy2shfv+Hj1nIJBXVtoYia4liQ
h4GxTe7cvvmaPl8pIR/g9s9vOaIKPcJ/O4AJKLD18oNjDMK49zIzAsv3W8c8IJH/amamMrp8qo3V
YNSnFk5TkY/6O5sG0fAePg0DpVX9YNrdEhehFESCKkvaKjmIY2NKUpydtqHYiTUk4MpkhDy4Xq+z
+wqwEi8k+C3It/gl3414Jl22Lgd6JUalfBnDcpPcRN72HkeTDIZ37b0fqQ02tBKz9Vpy05VCTwFp
FIawrUNrODiuEr2VFKaS6Yt4bR8sUWeFhB53+RmwWpyiKI78ukoluhu+/qQRqq5iyN6dgg/Dg/TZ
q5f9LyM/fnOfOH9PJQPADXGCUe4Y+60wDKkyMCVYFxb/hw3z4+B3XPxu+vJh9O0Odjhq+a5amGhz
m+lNnHac05RiTblGE7mAY49nVFNVxo7TzLA6MVIGwx1EUH8Ci8FCDnis2glY5fHRmxIqsukdSqNa
qZObfslnV4lZrd3CFtDDRtfkNe1nN2/Ey9y0OrFol9OQ71agnV+2UV+GMOJmSTdAkc5rXZFQGbQK
ZluIQ3rdVngM7sDfk+ZVvBzMZlMye1EG+NA18c4SnctqHS1UqoNYCVKe9pt+BZ9K6vNp7J9XqT7Z
KSDUdv5uoofV0/tCQv/ppkX1k5DuRrC3w+oQcxyWt4HUaWZjLaIzNO7aG6InJ8z2y76kmHwrLeM8
ctqsPCciGoi8WUnaD/Kg6KdGuQJGOy1DMsuyjB8cscW2PH1XHf5bAFhD47WksfrJdoj02PKuuIYZ
87J4Mt3O1FewHM5ZLglEK8onJOTyNa5LxJLfuR67bZTp09zwsKIHxl5mgwR3rg1SjqNhWjtfpqdY
9gspxMHB1bwoRpVP9ufTmhYOIbdqySamOjVBau9P4AMkN6NcW+HNpGFcU/4rZpp1B51Uq1Gxl6T7
J62ONYiMThtlBEPAcZqMAmx4yOBk5xxXLygf4DgJ0qQiG719ZO0kfRM4rrQjpzVK1wPHCjXDccMY
q8e4wIEL4l0gPPzbD3Nf/F87ALwiEElSg2B9PWx9vjD5hqjc6QUzNprRRy1+fNML3ZtVLIzjFjsJ
3KaIyuT5d6QAKNJO2R7z8Y0EEv/3P0qcAHQ1NTXbs8RhAwbXeEeccmJ7rqJOLjJ4gncDYipqb1Qb
MHbHr5YvmWrt3IIAtCCFSGOmYKBDbF55S6YJoJ4m9xjosIUo0gj9sIF2ZkY5U0RCkcTYEElo23Ks
OLw3z2jV6ol0ED8DmMiZCceFJI/K9bAwPV3JoZiho3GRt45C51cRBvO1Od2wDrOkOvtHUoYUMT0L
359n3d9Q67g4QF7BbWzrjt97iKTWKg27pBDN2V06wtHf6shHPfQXPDaGHY5skdQU9abz7wzfYKxF
3SsTY7FSAo/qcreuBtKB09wlmrlgg8m5EfjMf60lFiMH0Za+RV/+20lUz3zmV7fCjOCX7N5JY4/h
EyN9wCu23sctT19ZXNZsCg9CkJBvzrn0r8gMDb//0PC9YUhEvIJkvcmxy5QxtGRwBDCWySfBd69o
r2+cMd0jDmso14Rrc8DuNxeX0120Bq5vyyRVRlnT7F99eqJaWyi++eC+pEWXt+4enFRr+iYpaBQx
YKLdW7fcy8Ke9wnzntYH02lP5W9tZeoTvOH4FcHmay7tJ3V0D5uTs4fpwza8hnFVMzwBBihXGOYi
CA1IxDiobrnGx5Ppuu87h0wR7k809YDgE5kSon4+ywELojWOOja/BCnGTnWc1A4C10I+MlURcsvU
EqPlv2hHKwbCLKwd+mCjhZ94CEfEveCpju8bVRCn39foiKCpuO/g36NBIRYau7X6nila5LYAD0IF
iAAK7BaP3mkXaaXKUProwSEG+zuI4FdI5vje0Cz0HYhhsw1I1TsiYlbaFZeW2opQ9PcTly+ct9SB
IBLUSzphQWC2YbP0qXjzRnVpC73m5HFxjYIQiCByTtDSr7WINNdpo1iSS4fULLmgSjNm03tcFErM
tfU1+bvjamdiskQuRVLy7L5kYuDNzVwIwjOrVI+8uEfYENSp0+tk83gQ3nMes+kfxOG+EEKRmL3V
05xOIvEROpO7NLLN6KQwtWT4yo7u6G+HAoqvrixjffpmMY8AjYhKFY2Vt6OOHOEMRbsxLN7HB50n
e1WNvmJhyEVFjXESKfGshYuA1s6qkldWZscSStHwA3yy2aoOYHs6abPXQ8pRqEu+mwl4RKAR14mh
6WUgoFNhR4OfuYRx9zhKqPBinNJM00dld0iTDXXziJteoacw4mBWB+H0wib50erXVET5qXFwwf32
tem+pXcd7tfTAJ7+0aHcqamzrsdX+B/ZR3Ou1XRLzrPzJEcOo95t+PRMYY2YXLbrgz+X6RhM6ZC3
EcCrBlQQDNovhDgydwyt9QmL6YxzXZLZqLawxbP9rj6IKOaCVv6PS3zahhevXtFmAcUSuKaisCSI
AqK2JH7m54/Ox4qoEMT/vM6uiHfYIonpEqc2fX1or7+3+dQA+kJw/Cw0ctPZKZ/LE2s6b01tp8Su
8crpRaaU3SCeC7h/ebnZbNsAY/BlNw4ywflHO7gPXSXWrygbCexxhIaW6WPSXdLrDaW1siTRQIEY
7k3mmKELkMOOMwIV4CMs/64EpYRn3l826U0PDZFWn7m7uxHVfIg7E2VoQum7G6dHqi0DIcmCo39i
T+tdPczz1bm5KR5n8nIY9UbxbVgd81I3pe7MJz/z3syIJU7bSdobKMSmDkyfhJBRf3zXoupUPGO3
qWeEYk6o+ANFRBVEw/MGiAbTCPOPPkkpgPdOcruoStt7HXWtzmlWDvdJWaqwsocUIGgJiU6Rxm3U
dhYqgHyv+2eWp7Y8emnwcw3YQUC5VU9u5PvsJlJHFG6JzQjCBYUf2o7+1DKmsPUPiCVlm3vQFtDz
SJSu7lvOiEnOWMHZ+55PKLv2W21zoOTGqKm3pGKdI4eDw9Ao++2PfrvvT12FfSmHn8CVP7MSZ8uY
AogwSPvVfkOhPWYAbq7PfOkbwRy7YJGEkBJ5GmP5i0nxu9Hc1dMGYAS7wM/xTl1u35/ThDnNs4fO
KVHpmAUdpub2A3rlqmIyLL2AhET9JZZlifDSlMMoThynBI/+eIuzlrUjmZmaLxzFoKMgvpneynZh
HFc7hTNirsSyTdPPUBq+QcQuvOdOKcXlmWd0xbfvfoTc1KE+kuvYk4Phj6rLqaTOahD18BS+NsiQ
/w+E/XSpEBjQSD+yq3bPnqwBgxkxiEQHGkZ0uR7Fg4N3dfyT47BwHWYZ2qcVmW70SxNX+aZdEa+0
g+MVWSawRvmHE0iyy1wNyKPatWZaesFYQGDmBAyYhRE2uJoeTmhTnSioDG938Ssm7E5Q1zN1i+Ra
ox6jt8pLEXbx1Ahv8cSpM4CEB/fGbrSDh49TYUQqMGFhP4MgkVdKboqYi1pIkPVYzilci2Co771v
JMrWd8UhTf4IXYQf8+EKu7oR+jNmPmju9ylLCB1hhH0+UmzGhzRtyOTYK2gsnN90NwRQs9Kz91x1
o3/3QUBCdOmbiBDzXtX/K0jHLvVFLT0N2ji0KNXBHdWTMWXjSyNYF5866pYy7GXIBcTfZL2D8VIt
SSioHvpPdcnCiMq3CeUD7d5UHD1I4DI9ehkjYccotzO/+sCPTN5E6d1eNET1boZE9YHr+IaZtbVP
5nssGP6eFirsq3gwSKiK6HyzaWo8hdKYlWTXQ1zHo8hz7743rdGxvTtZcXN7qpysKvBdm4e3Ge8f
Rl5DCThj1Y7ri5jVgnuWzFgS5eem6qcsVgPmOhXV4AjNGMS0baTii6ttkIKq7fl4DfK1TQ+6hpNO
YJx8MoWIjsvUkbKKgzz+5kNJjbzuKfjwpKR189ag8QFCjI/jkmp0QEZfqxtddLlsPifQQP31cYpq
0qTSyqCVxUKSTXJJnqPuN+GxjMFnhkTuUwg7ufgEnN59JJDrAQhnm8E5tXlMA3k28523Ju9Bpk1v
7JYQh8sOFihBakquHhRdy+chtKVhovnFCtCDHJFaq7fBL5EDFL6QPb6AS00ycyG4IguB3MmHwF8c
s58Ptlo46JO7XhemwZd9asOoxVxy4OsmmjG6tl2Kl1GfiimP/wD8Tcx/cNtW2/m6iATBKADGxZRB
c+5d9+dFPwSTb0/0pn4YU6jiMkTUAqb5GjnBVSXBS0IFeIMS8i62wOSF7E0SGxzm8ilaiRrmNHD3
/GnxuNRQF/itpY9ThHbbfBLLO/egoP4Uc3enmvMQuDdOTIhwdvQ5XKbBkuIKvfnl5oDYLHOduPWU
KgNav2fQwB2+eM5Xc4H2MnA8ka1vlnwBi2ubW0bXn6zPae0mK5SYGU41kO58KKQH4BFEQ+wSgCav
LDXQbXC2SZTptPX+LPdKum05GWF+HCMqSw8L6M93SFl96ng71nJhHOceoKVQT+cXdzn/tO4jC7FR
PDknIhOtmzpa71el8bIvtxOf83nEbAj489TmK1rNOXTwGkpyNGDzGvb6qV+rR+Hno8caYI9oyb10
Xba5BIb7nOIjOrIcZXuPA1eXOtZBC2t+jqIZd5gbgTsSK3I2lTkpP9y51+qceYjZN2HwJfmSsGHL
hEwrrbL3id/JF3Dds3FzW+X+ikM8TDwCV1GrO4AqrJ4C6Ebkm/u/ix/Y75MAujTT6n0TruYLrN6T
iaKlYZqCR76p7WbllzqSORwrXZKhIyOjs3rwimXc4QqJPRKJvmVL7cpsVfrMj9j506FrHBjppgZ1
xIw6lshSE8Lofq2C+LxePdgoMlzl1Z5IBcyx8AAzP3qEA8XZMcVGuzkxbRTq+gAvuvD+33YG6Za4
RtH5eIDoZa1m2n9WVIEx/lFTfs4RJw3zbi31IAwwOUp9GNz9q9VMxPlad+CybGeHgzES7HDoKc+w
SaWNP14zM+0ligojtPQXiZrurIXg8dc8VgP2hIzELWFo/rHeEJ3ihG82cLYniJMq2P3t+7IQWy5L
/sfOLZ/QLUHSxyWAGGyrYdvyGgk4ZqKUKES14fJ6zCDEFOMaL+W9xJj6Xp5RdcZCcYojiGrubgVy
hs8+1/y56bPBe6iI/c0WJ83xemx5pM2RhifhCrPo8OSvrb2bS0BR3P2uCR4a479HfxOB74VG6wEj
OV42VScGXeyZneR0K2QoV3DvjztQyX0MfFI3SieXVLZFG5tPqPYk+LSl/4TDmtY7a7u48sYwZpnH
I6i6UjM4wSNZDDb6jMRsx/UooWT74cNixcPXY8Ne6/6WqwU7rlVqdTOaOF4RZ6m7wHUnnooDgkft
QJMGCvjHO8ffm95CksJeGk4q0z0HqH/SzbNi/cbzw7tVp19Uue2cgvICkCjmNyXr/EWpXByvtDD/
cGvFnf6K40nuPhTbUr3/4oHU185bnJ9CvZ0V4/1Rmh1rRnowlrpxXzOkJw7ggweX+AXVS7DWq7GL
0HIqdTto/BlCnSpub5Ifvw3bjeCT1n2+yKC+qGFOGf+mD6N4Iw+iVvMZolBiKpqwshm3sKmEQTlL
qD8JgTSqbCfgkOyXFnbMpYx5XVXD7ZxaUvQ6gHYz7r0468vk+d0qktKNktqXwL2xV8bHV1YAcdGQ
byeohJivpnc2RTu+4L5BqD/GNO49BvtjlqHVbmkxemU45MfAPTQEOfttha/bk+p2gm7xAfVgrq3s
2sKni8J7RRPgl+sp2FcELZ38VNBRm4IIT4gec6U8LAvUZZuzKjg4mkuB4oWL4j5sSS69eTLkKo6R
f1wAALgVRArbU3gpZRV4SJRgeCtPPZ/exYhyRkyeq8PFxShW6vstfm2oUEQW+0q537FMKCsXZldo
RlEGeMf7Icg/an5aXkZF8CIp8OhC1699ZDMTEboQvNfUXFCg4BKaxISJ+2pP5Q2PIebVuQFkcSbr
U7kKVRQQ7cQfCvOL9cMIk/qD6Kr1kxIjckvHfJuO4Jp8tr0iXrizUBongxIVky5OIZhhPkOURspM
jZM6+7u87w9h1wPzFaVjVoITl2JUxN8LYEZ7thPtZ3muHWaDbo9RJziuUwpNtJpgBNktRWTI6f0j
cC3yKWqj4BQ85A4RI5rC5erS29qYHt3GZZz8tNf2qsoSdR60mQDV5D6JyJUJRcQ6pwmrXm8z7dfr
Qd0iFEHBnBVwZC8FJoYjibpNdHxuaKSIBnzpKQoInlLu5OIp2923wdog3ne4ZH6uul+i2ZjWIDEw
1tPHLaqcIR3TV6uUeICYQINUQ5L7o+aZZZRxHt7kJ4m4uMdef6elz7RhL2ZB3co8D0Gj7GJK/HCR
is3Kqc+cfsjuA2vwRaT6R5D3xJ77ISfSwPT0x5rwHTsOSUfHR7pou8AsMxUYZBS9TkfAajm5N0L+
C2duFIXfawHqkrlzHP1R1MmEOijP9jDCXDCcJqUTLSQ3vTOdOuNJB7NwY1e9Ohg1PkCCXWeTyrTh
cTghvo4zMPLMlwORsNBOr7rTwcf2Gp+gIcxhJAxiqYkU2RU3hdE7oosNLv71x5GxCg/wZYTigzBl
aUaPpLXovPEa3L57H9h02f7Zih7KqF0UnEg26y2UPh2G6OzqaxQ2aOrzRB4opI2hQwZ6GdVyFd2T
08o6t4tYs8aKXVWT5JPoT6JBD8caaRt9JfODUCp/pd5E04gdh9FJTdo7hvTaps6Su5OpobDZ6lXf
JWtlNNqwA+Bk3esyC5GyJRjxKEUgq6xpcTN4lDbdHmB/BA5JJu+ja5ObHtEozvBH4K7EkEYMUs7d
ZKezX4aFen9E9yvS9SIJVjDGr2bo56fRFZG7HrMuG7ijN7xXG9zE6k5lEOx7de8NzoNe+2QbQ/KE
E3X5/O8qMo1cD+X1GihQ3RqP8fHBA8NJ8kpKy0b/hQ8xQENQbcGaWUAkOqH69YZMz9ZuQ/q8REjS
tMKHHdo6OhY9PBguoxW3kjhRSmBhdOYA7DrtqaIWOZBabNuRFlQ/1PYJzaxEtw+m2a69sAa+GrQ+
9Pzg156IHodHMUkIxtonK9Hgf2H+UxiEWETK5BeDg0Lpm7FMNBn7bkAt07hDPP7Lhy2keONN36ii
66kTB5KX/V15SI9EGXDTzXOwNjwrWCYdRcfY9BsNMjvPJQt2oNfhcsh7xJX2dthO9w8KWhYZG8Ly
atAczNdTeKSpkBnkFmqVlol9hxj3xUfZSIhMDJDbgxCdbmC5Epp/YqR9SgcDkR3Dn9P1KwNqYQfX
i/6+HkIM+mURy0Lw5OeoG50R2Tuhdo3438ip0VrKOi9bMcR2E+zYdprdFF0zooVUaQqeOApTM0fv
GCSqIXcUTWdE2w5+MInQ4DObjfq8gABu++DnCLxjJfK7BPsqM0skKHPeZ2wIQ0iYQQd2D0g+hWRm
e4NrR+JFeXcTvRHnAtA3/gFeYAVBz1rHRAvEfn13IybVqLyACn9yPfvyv2bC3Cr1F6xP/vGYM26A
v4R4mklBe+AHM8RpATsCigQut+/01nKkL9k54BSLvSV41/ZaoqvYKIuQcvD0zegVF0peZBGSQTpM
uotdFvAGTf7tZCgq9P+bysk5Eemm0uGRExEHGNZXoLJL6cgERxmGTVIGsauWmxDFy/ZM0Gf0lsfO
fbXa5hBRtmjbt8g23+Rq2o40S7ya3VDDd/hOEkP/BJ9+YI20+3jYG3SlpIswWxtJmPPAh53BezWo
WzwtTaBS8sNK4tm/tjoeU2FpLLulIUORb/WonmYxqBEdCdPCww2cfzp9mgBdLG4yyhu0GkGBN/Lz
9Z3SNtAbVkU3DmZo5CdlGDjTg07jgfhDXZZbrN0MRsIsaoxhMkGmOlmkDFLtU+EuFcMsR1jD6YPW
N61F5XDAFD4LIK32jAlaeK4xbgQGMitmJb/3R5PQlXmqU18aWTOAvgl0ebwlx43vN8UW08dsr/oO
xZr7pY8VdMG8ArOU8qnha7L6pPywGqIjXcPCtz2f2svfMfvo4we+SlicM0J8ocOrCewLB+FkOBcZ
+DlMMpUuSseKsDq92b3fGCBFjnP+iAw0lhSQFDxkZDMixleSPAvqi4OE/9U8dLGgrYSX5c/TUr92
9iErYllie0vGiVOe6eEPPmmay/1NM72aUspIbBu+skK5km0tb2gpD+kBKpOGYKq5Imtq8MG1pFJx
eQCv1dI20XQLbm2X7j2/vl2cNHrqDUE52WtjLfFlxexRZhO2lMOL8W6kSn5YVUB4yqWBcaaWGLZ1
eUWe48hS2nXFmJ06YVGjAwQGeWs4KVVlSOC88oRUhiB9pgsF5BaBlGrHi4W7COI9XW1k2x8wMxEr
BOztIxWM9gP9DIPGQrhTaeklz3onr0J79/15rp4xq8KpqyRSPkOQWreVk1FqCxYsx4CyFT+RqWKe
RsD0j30R/eFQdUxJWaPOin7ImTLWLbiSFyQecmXiFA+KHXLP2dH6pqejFVVLKNgk5sK6jcj/T6YW
dbadRZh4tThT5nc9omgw0C1m/dGbkfwndrJRbvw6VJOsuSV8Eh+gQ5JjDO/Qq7Vv463xeS5ODtij
dOlIx0SKEnbh1MSbe7kvSqelT40DEmFThaDbkyDZuBmNCBtramo6Bm9Z31HreiDfOF4GRVu08Hbp
4kxNpY4BDis+Qf2YL0Bns//+vbtaK//Uy+nfAW+LhxgolHt+0l2hJ5mPf9s4ppeR8b7lq5t7/jsB
aQlAzWo+Co0YcsxijbAFPdZJbovfNWLY4ITa1annm9mBI3YuGPtYQb3JxP5lXK2VrVNEdvPG5u1o
hlB7tkFPaOMsAEfuNdKkd/zvjl5UGON4ZEVs50h8de/pCHurw7MY1L/mkEg33kmFudaMePEQx0dD
3N5iol1DEI6GBPzCjfPX31K9bzvYhuorexaUC9wXh8itB7vQmrvmVdwRw/spZ073O2W8uaO68fZa
UF5kcm5lmNPdEaclLRHLQD5xn8dMPCmgorOaJVtr2pQGRHPbrFnZUrx/dJ5MxsMpxvGexNtCo+Q1
rpIFU9k4+gksNA7MkVV6XiV0/FABRG8rKPf+0ZppNu3jdaR3CJqZ09lXA9pX0OADPIeH0nUOxWa5
Om+7O6Cc25ZqX4/HM6Mdc3gwIbERuI260H5nBV8B9ZNnE0M/w6yexcshfgPHru2Gdks9/YZyt7Mo
aRKu+ywJsoM+LxrDuE8WOkC6FbDjZlNJRAnm8XruZFvLIlM+OZ2C9MIGWtjoQ4qrpQWTAE4JZa4k
2+2dBt0bXbZWs3wU3GkoD5/GRyOqiaaW9/91/IhAy+zN9TU1kXnHbdPLdn6zcNLt4YLs4x7QeOSm
11bl2vFlo5oXfUkXj87eIfXPeftV1DddYRWuVoWyGNq1s1cGfRe2fhzx0f4YwPawqvshB+jxPe2E
zJTAdjZ0CpH9G9YH9iPFNugcS4qoGMGsglDWiSn1tN2o1W27cFonU2Y9Qyo1FmJuItfEdougU48T
1QKox0X5ln9P7hoTy84RBTlZbjM3v3uytjCWODde2/+IL4qItlq+yxgKyp6n9Wzs3Htmbv2KmO5F
d+JukzCWgibi+QBjWWQEtRrfn8aWHF1O9lbDO39i9WbRzLM1GZRDYkj1t4S9l2WVNgZiiP422tkz
cgC7+u7b/jjAIi5KP8zrNjVpXFnfCpzHYnFpV5a5Y9QEC1aooq/WSyaYQ/84XuvDG21krdsvi1qG
WZNreBYPDOa44hlvfCJlPz+XlB/XzECZHjXasvVI0OXBprmS/IS8ccEBjYuESX9LUyjNPYMvoH5e
GHaVHnLloL2tfCsO/VUaRBLnd2zKAYx/0tSpRVsB9+Kaer2YmOQP/a1XjTl2/WfWv7vZlACbBY/j
OdtA59+XUwL6fNoOgVqwLxtW7x577avK0TEwCXTFJgGGy5wU1GNLWRW45Yi+BYSwjIJnLpZaEbSC
CNB/hyU9piZ+dKT8hPKyBosdv2Q2qjLbeNa3r83Ie6TRg0qnU1ntm7VGgmygmZD1CP6QjNWkCk53
/GDV3pWq7CE4hGy9SqrBe2ugR5HWN3vBC0mUitbeGkGs1wAHlcoQvVXl0f0t95s8mHAhcFzz2X3f
FlLLlDAKqgTFvYNFcD5e6/flH4ZXVA2hPMyJHthc8O8+Ca3K44fNUxJfz05DIT5Y1+eUQ7lDJmPm
8v0GWKfuiiT9KHH2M+wy6pJ2XlLGxiflfa0R2xeRdKEEluFKSltPk21Sj/KozMIEF5Henrjc06vD
0UGPTbFCLDms1L/XYG1K4lZ9lNZIwIb9o2vs/IipebqqJTq8GzMqwUCn0mzWuaDPgRtKMATsPjct
2yZiCAK8dGo27rvbmnsAGRPAb+wkujh3Xk2HSjl/bo0MGv0EFV+W3kkZeymW79aBbljEeSEtbtWu
dus0MtnpXpQDFFtEZvAfUI38a+vwjJ//uQYbxEyREuosb69gOITRaJkObF70GHte3Uuv+NksngE+
O8vXxZs2Z/xwYIgNAWI8KStzlX8Kg4/Q3K0kOM8819s1hkdIet0FxrUqOXesd9qqQ8g+0iY3iRgm
ppJywiLRSViS76udz3EcreAphg874SnS8MqqA2EhCIYYAecv++JlAu2F8MILgGyi7RUTh8O8Z/mP
CN0JPvmjH/Fk33UaX76/mdA1ER4QH0/Z1VxEAw321vp4qUswlmIxQT0jsIqgGVs1s59JikKlKQ7b
mvx4Tg7LbxD0d6MlVPDoX2vH4REVV2bFnX7TQOSIVVoWumZd5/pIha4Ht40xDgI9ygRvTgfYtIQC
wdBqmvQYXixt4g+SKZ3nuC2e2/nqo/wyYYDYEi85Nww7dB0K/VxLPdW6e8J61M1SRaAPKt2Vc9tW
bmE8X5wkeR7omPl6hZqu9dyJZ2RWpc1ejTsoqLZWoUmBaqEfhP6pHxvhmlb24qGQmbDS4zOX604N
K2xO9zg6VZ0Z6Hmd2hdWmSnmLBU3aZf1RVRiQFvgSuuz5pO7A9pTT9AU7Y9GB5+5D+bAj9czCQqy
0IGTOKScab/PBitwDGqdkDok/+aiunW2UHJA+svluppQmb4OuXXXz9u8ld+XBJLnvP6ZlGmuQLEm
ugcp1BPnFaxva3VdA4m8HiIEiEGvwW5DR3wke6tuY3oLKY0TvhCtIFBpcRr2wCGc+j1YpAUjw9AO
/VVD1c/WBNRD1OBhQye0hFx8FNxsf93pGU3CBxavmeLrBxKQbBrT0BzhAkreXEgSA8Nmfc+0mRSZ
FILYE2okA4uQdsBfXn0oxh6WpCkPjq8wVG/QDPbFvHEY18eDJaA/UbOTXzUoshrJDCp1Zx8lu2R4
ou5Z2cSXT3Tb/DR7sGQ7hDFcuu+tKnDrG9bSlXLRxZcz2KVW0OQnmOci2ctK7PKXxysUu1/0D9Or
ehtJrQ0X8MraAJu27k1qdwsN2C+A9RKTk9KHyM5V7BSXSiPRpRjbFmbZzXP5Z5HAmh30qSnYnnhZ
xbq/n0bIZRmYCfy0oj2ulAxingdOngiEmQLB2m97YLxYIcfEVJp3Zz8nKLpQ6sPcnqOvRT0D91XD
KOwgendEO68MgGCpUG6FrWbuGcQtOCYQqwu6+R5TB2JzlpPi5jZXFfHrRZHmXp70URW4zfOCBuWK
YrM+es+YuGFERdn/kn5K2lKJospSqSNReBH9ngTEzb+iumOUgTc4VQyHK5btVQs/DFxwq1+1hHAa
U+y1Wm/JDwGVcHYx6rtKCnC0j6VMURQhGw/rsZH8w84I8jWK2jWGse4Gj1NwrDfFAZkSqDe4Pf+1
l403ujRlZxSv7v6onb11kPYjLwSvohO85pltkwcBtLiiN27zCrCppRxg5QqV/0jh9TdkCQ8X3LOd
14MMi9COF7dxSoNfsEL/bFsElvb4fn6bOJrw5wF86yhROObFNxUxNvPKcIPrO5tZg54cUH+uZtgZ
Ay51uX92NmDV+cKF5Axys6ww97jS8nbetrNeG8WfaKx4Vmbzc2wUXcmKwEq4o6kixdfwsSJ//Wlj
euIfMTowWHvJAw+INh1mhYruoehrmIQPbpAmwqJ6kISuuO70+IYozIt4J4pu7WzJw/P+sxalXksK
wi1RH3Tn8P6tSSYZPz6otJAcH87SIaaaDb1ecBlfLpeDvSgJ8kHoGrsHdfchxWXwiq47bPpxFCGf
hZKHkD+JTG7UqYD1RSfTNxkQNMkKm7S0tZPuOv/qO8HQ+gbtT4vFvhJRIRWpl/lJTH+OKHq4XQIE
++LBvg6KBl2REh7D770aLmRrzEv3MuSDZiha9kOm76d4KI8g4jocY5ScGiv0u6iEP1aXNT+361Tt
A0EGm0UfyKSpdwqptZRYqWerCzbib5LcfkYIrmQ/9YpsnL9YYWHDeWHeenvnxFRa2ctRDy13X75l
NEy8yAaxt2ITlUHqZ8qHpp/LvNJjTv2+m9HyWAzc2FdFAh+D4YVf/9uEGlCsdJKH7GSEHiAqaC+2
2saa+s+iKVNZs745QKBsnruHk8MfUt3rdWfBlyvyjuzDo3eMWZ9SfsapcJOln6j5BwF12iW0Qsza
18uZtxnOoYIUskGqBXIqDMlO/Z8VGH3VlwdCM/DpDPOAMLH9BApjdfaLbVedXpemDpvP5PRGmJrG
W9zYk129fiATQKoEdIC8oy3c367XJYYLqbcdsUAZ/wQXqmaddg8VO6aM3znLji2W3Z9XVkSHPwC7
J9NMovnODvJuA5X5YXtcYDB2gDnMBzr+JSQwk7fY7ba2rzf7PSJatsUYi2BueJhYlTH5R9f1++x0
LEZXBhPEQpfE2Uq6UkySMqQIPJPXRMxxXW3Q9K25INkF+vm4LCJkFO6dTzRJnY0cjG/fE6ClUd8d
pyQvT0D3T1LLqN+yWyUyFVC03wheKBGpTUQ/ayRXyjSUrzadRPbAXOSU1nJu1D4XzZRou+UzjlCe
DgvTI9rEAhNmhZ4363Q9BizBjjUcM+rT8s2uboK+1BhW+8qosKbI5IZZnmIJqsz1WDgfSuJXXLaR
IOASOIy0LYzI8FcrQwlkXLutWnPgAA511MajffTlEWhcnElXzjOylDAZAaO0cfs1E8ZLj1VfniQw
RWMP1X0bR9GEeSMB6S7QMnZW18fTO4R/Y7w4+VgGvvZ4H3SV5ntRxXIaaazbiSsSNYj/UOsps+9s
TAYoVTGFOJ74VbAokTBV+8aFNn8Sap+uLRsQa0ZdAL0COiSBQLCIdFq7qoa9clAeAVREQKshO/Iq
irOWR+Dp/C5HONRbupve55gVqNCoQl0NgWjE3aBu1Oiv0jUVC6a7+mq+q5k098Ixca4Mrm5gUxB4
TM9rw+sJdopgZIzT++kAyF6mqQjqkGFD5XkbVtA+bJg/WfSyOVcjgrH95A7pYJ/UvtmF2axQssQ4
QagNyuXfpw6kZ36yWxmwyRt6GFPKkpU4sHxkOEpUCjmhpwL5PTJxug65MmNfrqW3XVWjJKh3SnnE
APvG5tdr32JObkZUqLGrp8cQZDed9rqRfnqyPqIFXD96ijR4s8LqoyzNUFde0PRNKMjKLssCWwuE
pL6PIr3LbMmOSKuclQ1ICH/vlNC2wc5Foh42aiJmLXKJPa9e9P9kkzeYhVQWJN2MdmTWiFtOf5B3
Kw+uQWvjVNx6toDvoY8c+5g+kBmvcrnGRMwdVcUBLYAiTl5FfKZTS8HngwKQONwdx40q6RG7qMjx
Q/0QwH63QrDiMueVIX7FQYYw3lXEuNk3k8EIrEMHbmo8VRID0vIr/H7g+p50stofoaaytoFZ490g
iw0L2fdGvr3QiXtc34e/h0BpgGPMeOsBAcpA2YnkmPFu3PfmyJJoW+7l3NxTLDkptbcGy1NPcYXJ
SHyV+cWqGtsELv16L8n4xBNMxXx1yaUVVni4oj6Ud1dDf+Ze7c5yhoUga2i67kxB5vhjetDzL7Iq
O1yjWFvL9/vY0SRVBN4hZjKCjxizEh5gFTN1sXOXySeseJbJJEWZIQbJJNrrBuhuzeNFQ01UsYRk
brw6O7MZJqiEhtFUdWUS+ZwNFEqTUU9AXyJYMQxj8+s0KJD2FB7975n97VZu/vhUSJvdid/ef9CE
w+Ee4ce+MU/g4QioxSW/5D9gNA4lRG7t0Cjfmrk7HUhmtOzP6t+xnFsQ49sP5WXbZqF2jJoBlnex
5ZXVLNgH0gNhbB/S+lIeSNUPyiFW2jvodmeT+Lwuf4UTfCoylOez66vq0edBXu5y1S+mvI03Fbs2
n0414E5FReyALFmINEAfMfrRGSvn2pk44npFwzVed/9G36lIpqehM9o5i/ZGB3LxxfqcpKtiO8+5
gbyETIOtqoGqq7IJ/7xOB5BtPkNl6txHKCqeJQdiRBY5ct3g56AGrfHIvNYB9uDRGJVE/cvGPJ5U
JEcbk8lAAGbe5IesOPv3E+ocEHqv3YONBckEpSJrjAtc9DiL5riczosmCRtZ5mLmvENQnkbvDw5q
J9PKrY8tQy7Dxkea7pGl0tdzWfJhzTlUFlK+RL5UKoKAetMeNhmzOVD3vtT4+KJkuX44QpiPajIt
/E++4uNb2HVnx0VOjIOrIOoGk+hI3UWk8TZn8WZlPy05K5scMLLAXh2dGFd0m+dy/buwllqZHSls
pr0vKtLXzgcQtZ0mpgsuT4fbJXjmCIl5G0PVAqDkstR6gOxCFcJfw75AfDvqlv17pWJx5wzTol+6
YaSBV/hcp61FSmbnDA/z7rJfLyksUh/WMqUL6pv8Sy7f3CagoEn/pDCc9QucktyMSYLNFKpCcYAC
9qupJ/rDuB0n8kDq2JMp/YgvHUUK+isiBgSgXhUiBW2VykF7LAQqtiD+oYkVtTo3vqmCi03IU/oZ
Q0d2d2JBBXYUnPCr4XFn7NP1T9dvPeReMuRpNf3tw94DfWNS8VxN3eEgQozc7qi0myj7X/6xcRuM
9hf1jraYdfsvlZaoaKMlOPWvghkuHc9sCYVy5Lh7K+RaIOqpCa0KB8hwwp8PFQHxf5caNjpdIT11
vpo0F/0rPoJDu5YbVD6SVlrIiqON9dMum8kS8ZZGg+s5fA2oAAUaId/v+uecUccukA4mPI/DUMh/
OG+lUmkdcC158Yfc2YNe3I/2BGYOtGw8UE+h1APHyrPDeorT1Agnr5u14NF5b06xJ68zvuzw0gsD
MUhfNcsqRb9+RFYWPerCNd80h38CFN5R0eYOLdVqrV/kX4QhnyRyJsqUXJQuXTFMW5uSmVcQL7qj
tfUkBg9azwdhsVEuvpoZRwt/44E+Q5qROUXvWcUF+d6BD18zjecokUiggNI5BxL7J3urEZjQLQKv
Xw8K8LpQQ14H4QPJNZIspd2QrsSmKTuTKbQtt3p1q18n9UsGNMfi3nY1qBzq5JGX6Tkd04T22BDH
yfvypZtC8qQpKu/zfTq8mPzLMa6QRWQ4ZNazkX9i2wNtbcEhLTe3ZjMmRViwyPkxkxuNqsxJdpAt
yPTlu9UUJXRNWVA64wMw0u3F08R4VRPW6qS+eWUtbPPoMTqceMKBvViRPff4p49SXxKzGkpAeB6C
rbeS2A0K6CxhU93qwh5gyQT1Fw5vQK2O9syw8pH4KDx1BjAb53MGOrPdup+62u/lZmK53rEKFPS8
HJHKFdqJYcZjuBPNBG956oIt6sCQN9Q4e2/38Sm3DjG+KHUCoLp9IYMyeNeYvyG5y7qIDqdS0znj
4CTIZjT2upinI1YednkSsmcW1eNAjaOwovEpzEcV+p6kodHFOwhGy8yJqfu4XAGTzjIF94aaZdXC
5P7FlfkJHql26LvREF+ssWR9ugOOI972EHHnV9FkcCItX/abof1c5mkcGU1/mNjlgc+6m/NDf2fh
HkjT7V5BIsEy1Du+h979cA6CiyFW/ZQmPT1abUKf92GsW7jsJvkjLb2WQyKzs4aZpMHTjIq8QmaC
lVm7ekmkiaJSfL1+tY4C7GyOLIz/pltdnd95w99y27fA/bCXxYjHjQZtbnnm3uZfQlvEHoTWw99Z
LGTvTEmt/UXBiZEghXMHXQ3GMmF+ZTMuozEJxt1kvmvmjWdq6PdPXDClr3X3FO8Vf1GjArdwDHaF
h4wVYEOUGpBQl+HvKZF9WnThq/dKlnloWKOoB4Nb8ZO0ihUUvt95bzr+qR0879z6pyezrzfwXY/6
a0GW8JnafTVoNLvvXuhXwfozwWEX6UOLn8Uk6FtM4LbtEA3SGZp/F5IRrHk4sBwM8QaCGP7joAwS
/eOlA8YH9ol3nN6LOIEk6kwJX0KEnUW5ZgaMfMXn0cfwqM4m3F+py7OElyB/lRR6dQMySPEvtgZX
S1LtRTpWyTLzpZvCKjk6cH2NPnOffsgTn62PMKzMCmDl6S+j+PoNc8nQnGanWSll68W6y8ytm7nM
yqPCuN6Dz9MCl1gvT5cB25Rma8Tmmwp9W8xn4c335nxEJAY7B4iv94lQhY5K6Tr2wfA0W7o4YlZy
ox6uqCfusVZbJRYeg2hiH2igza22UIpC/g/TQMwFC70oxuTH6LPGXJdzVmR5QBY63flPgC+rBdxy
Fn2+1QGBKBaaJshUIQ5Z0LPeZFvCzHxRkE/UPUCfTQn1XZi8nwAkmIz3dNKBZpdMUAeUEW4qivPM
pLTjkEyZIsX2Tfkts7lVCbCLSr+TSJ3ydUK0QKZHEJC07ZiZ1wQG3oR9wDqyzhU/dcUtF1oRkYAa
mF8aBzH0kW0bKDSEU8o045R+od+XBBAz8n36zft2WSMAGuiQY1CB8EMIEK+jC3YNc9qRDN6tYaoI
ePmeij+wBJXh/6VtYQjgHUMxG7Rf0SQrLJHass70ahq8pVDDc5V2sahuaMrRKViEflmvPJS1dFk1
3EucDO1yWCbIZP4a9gGp29lGf9B+g1IT6577tsezJTNdVtBhpcGoM37f152MExwRozLjG6lW2eK8
tyns+CU9ondppdFsjN9jTnJC4CvFctdxqCQkcAn/g2N/3BFtU3EBlasVP1p1IioRE2mSK39xKb81
N7QJbnrHOjCeni1gvclOOssEbDPhHrCTPBOuyHfgUm9n+mXFfB5mDtaMuxedFXR0LejEbfZRl2ix
ZthN5yjW6/I41/xzMbgx1Wzx2OBqP6fHxn87gKDM4gwmfzF+3Hnu9/Eq5sGr0R3FqYKFSzG25YBf
nbMWWEg58bczDVSG2BbTE62S6bATHdAg4NXRiOincha09nHzJX7aEaXJbiqsB7fk7bNHAHUlKu/f
Xi7VV1VDoLvrBhTnwm+nuXAXMXi84N1tl5Xmdua0ZAEvsxiIj9rDSeqz41N6fuW9ef8t1W9z662U
9XFu8n2wYNZ3GcfT/xvV+2dulPxD+P5Ote/895kMtIGxXOp8NoAGvWWVlGxFCFWXr/hZvmfrp8up
aw/gLEZucv801x76CN0IFghNi2RG+Y9AIfZxQAkCoONB9LMmxBg+03Z+PV999X6HdrBl52OWKo9i
MgJuyktD4zoeGgl/iGHMAyjqEzUZOiTMpplWTfO/XuGXASNOMZrtGtlIznIFkL7UBwYW2KgUBMq2
8MtIXrXc7C9L1x2Pv8eliQYIjVJx9LCFZrb5KYi4PWYtsv0cx5o8xAlL+ohMUlBBzRbmS09aKDnr
tPrDdZ5n/0Ybih7NtzhwznClgScSMK8L5b6QDqUw90upINW/E+b5B0qwJHqha/VWCHW9759GQgvb
GZJTze4iBSmCjeJkts+b9LRqu2vnYFdeb6GHQP9zz4TQak6ytLQfqT2GtewHAWRSIGL0gyqDGSHV
tjjqOtud28jSJ0zP8znIiiQiS7JB775KjLLumdxe1Rxs2dqIQzD6JOh10Q+XILlXJDw9eSn6YmO+
0qXsrjJRIGPqFCsgFKJTfhlGxgkVZN/xdUNM36x2mSmwM4i6lv7A1RnpYrZLDuiUfpU8trTh+QpG
o1HYt3PWeedOrWGkqYv2tAHDA+oD4pxtSLDo9ANS9EvG8gfi4CbuYpghWSlHs8NDN87QO5Oe+fXz
lAz4Yf3ADFDVCUGc+YVU1evVBzqpGWYmYT/3hJ6TIjEOZpPtUFGcJrk7UAVVmy7MxYjCbux4mAh/
VCq13QDi3/V2yDXz266xsdcinE+zXreR6D4kqmDXuEqB1mJNU15nPy/jfw/CZjZO+jW556QMRVne
HcrvjHu/x+vOyH7QSX6cU4cn1H9/DStxFKCM2VJVRhKbfuOK3HHMTxit+q04L8nZH90bFM4qa3an
KtH254IkDvmWaQfqMxHvekeSeu5eBBwizkJz99blOc2J4vmWiWt4wnvN1wlgbbDOO8gh+RgB7UDq
/HrH9bwtWcBPVANsqmkVsyxkQ8WKuzunDsQFKzrhwK9G+/gmRq+dwWZzpkQZSsTfgHmyB57Xsdbe
Gy89CWs2PHZTZ9bEueBgbW5cXzdaVcvkWzYzl91rmZXzBC4l9WkvK/sMN83cD2WeDVQO0jjOrZXT
+rJ1llme6+hhtDB4KSgigVYY8NG0kEaaYc3rNDDiL/e+p46uuDk6I0Ylckq8uE8l3pWBOB3LbGZF
dvCREtxKLPCHbZonV/TtoJSCaA6/TIUrq9S3yZh2l0u7e5VFXfUv545KZPwb7t/WZpqCCFSrVErD
3E4yYxRf7Twwzh7gmmeK6+m6UXkTmOsxWGPs9NmEuN8npaOjfoDS3B+z+yD2ivfVwxX++PvHwlqN
Du50lunkgeCrn1qV2W2gvmIqsKAJcqBW4hMQHIKfxY/urivRlz/Zw8pmTk1oz1qMskeW8w5m3Ifm
mZmG5XHMZD3DA1fIFIhQUBjr2NzFhVFNjsCHbBK1gTund8CDOCwzIE7dYluNCR3P12x6zs2HbET3
5xJMUj4RqECAavl5bt2j9Lyvp8v3ufSJNkBXVW57ZxF1vgQjr5zUmHja2clq6q4q5OPbr7FLuDXL
EgVUKeCHLKlSG5ebPOxSRLnWJHaOq4TgE9EhCQVveR+fN/xFjjM9KQzE0cowK//yYpQiDGHJYodr
Iq1cOZY67uQyUNVXfG1qrxYceHK+WvOEUfWcEKhK+7d22H7zQ3PpsNPLQD4xK/w7gl82/RPJDkQI
TRtcWpLb1SUIvRh74dNUQ7uhYb4ISBUANe/rIxGzwXEmO6rZ+YhNqvX+94tlcZJkxnM+uvR/X7kl
CDGhHYJp5op4aIom+KS0u8Hc7oh+denP8bOjBu/WMsT2j7lZ9nbgVlmHRDx7chF6H9Cg+SyB/o8v
zHrHu7QVhgElamTsDGOs1nuKcbNYsRFbEMoxeAgx51VKA9JMdVr+DuE88E2GNux0gq6kJRf2hfZe
8PeDVOlGSU/v+ve+PstlQI+AXuKVhhhP1JZUhPHUihjPcH2tpfsyZ0mbzingUHN1oCNfdZXpXrTr
VFzt4anH3WntOowREtCd6DLHXd4ikjOKWgdLrSLlr2wBN/KsTVFHiiPb0dk7n00s4LB6/OKVb89v
+pcQFTSnFiD0duBrUW5BVpdhbjpA2Eil8exmPBlxtTREvcMnLTogbKZeE3Dh2SUib5XTJzHpxAkw
r447uMRQN945PHxxndYy+C6ScRPa+CHtJQiTbH/2JrGvUV4dqWO0Bckl5BX324HKtVlTQJldPEvN
XInd0kI1oy+B20+oAmK2qiHtBNSeJInaOnU+lySt8c31RAgwutXm7K2t9yL9CSk0ABK04qHCe914
L6Y7gK7BtCGwRnZi65mNgpMwvYTNKXQRYB0PtAuiMyHTiWmhVat4/5RXJ/8kqvz3dTA9Ybw+J/al
U69EMHWCfkELurbK3GQ2RPYzFJ0m6bCnFPyuv6P+iX788Hm847ByP5y7OEtz9CkJxxTav+xHoRMb
QGQh8Ri3w31uV5Mzsq4vJJfEglECWVCOAYY5d2Gg4A11K1M4cPGpEOkrjEFL/E6kukiDZfkgVNQQ
nIZSZFS35sDn6V3y/vKHDBu7PXZL2cFqnm9U2cS/AMg7YW0w92QRrIbSZu/QQDSMZpjmbVp8walh
c1hRxbQmXo/V+d7KtrJllzVe3IrBNRM3jDKpm/Gw3ygeoo/ZbHcfOX8ZB5APqFFs4SUMQPhgdjAY
wJnl6PbjBs5IjMSQRT5HGxp6JW+DT0qMRxL08wJP6+6m+9MpNZZXmt9rz3M17hKt9o1L0qXjYhZN
kjWFgPgAAFJSmfZVUjuGWzRLyFoXnyDF0XMDqTbAGDI5acumS1OGQ/JMCJA7oMjEAtgB/gmgpHp8
L0A0jd5nFBqAv9/14sMgsA995Vx25Pu2/ZCkWUMVIlyVoJ8xQAIo5IST+ZpUxFwr07PL0TjMU35V
g1OM+YbqOTZRS4AM+dRR1nY6fB7m1EN6nKCVhKfgF3VUNK87Y7abLLBHWPTI5rBnjIT7yovoX3OM
ssddJD98vmoD2Uy6L7rkQHEJlnU1NYC/EDzL1hECm6rl2HWmgli99xB7qVSW2tnBUTNGSRSPAzMt
tHc6Cu6qnfdP9DZXJJ2HfrotLapMidXuAlMtKVqXQ0Jvwnfz9cz2xGGuNgbRdw0IzH8rVPrhQsAP
iYSjqI7GxgkwSIkAPypyS9ei8htGheYb2bBs+hxWoDTxAYmDjZ7+RGGyYS5xLL5fNcih+ED7ueR+
1seQUw9W8Yg/w9ma/JNTfykhjxim8JNJ7RKO5ARJTUbrnqLRqJcnaku8r3Re+zIsQEKmkLWPlSgl
heuDmWFRxbieRNvVwNMYfQUQ1OyrCRYbsrc9KIfGpKf58rvh2AIfBTCBuLA+dL8J6bBCrDYYHRJ0
MK+LxUoHpB3UD6DdZbOtE8Gv0eJVctO9vjcDklZ0GRFZpJ/9YzNGnKM0csqmU8dVJ1lkR7pwPTcs
IGWCdd9Zp2UDTDR9QJTZT1s7/EqM+yAN7SLUhwbzoTyguAgnZz+n6Q31DC3pZD2ivvSbdm0REQwz
vaTonScjBi00lI7ziVPG06GO4k3P/xjWlxEXFLX8oquwsGJJ0oexbb01vkpbpCJAGAjdus7wmqjx
J4GTAs/AA72erTLWjMkJWrTX73BjbdZ8irn9Sl5fuDP/cp9DpQCahiEN52vzqzAhlsnKH3W//WY3
IwCn1IMo3Avmw0AYdK3HiZfJK5VT5ICSni0fp/JeEqh1/yv2fCOTH7ElmmMug8K0hprjyBIQSwXv
Ad/Sh0aNoBg31fiwhkdFWF5+Lbg3xnkHyItkyGtBFVkJiXr5UPYJk+aDTfGQm9wwWikNiuGBrCbs
GP4zZuEOkrW0Cth5ZdvdX+LW8iY0ydIVg2Y6hrBfi2VmJWxp0NApGDJjRHmVowsU3wJuFmJsFpZf
EqQAwNKlqB6KAMqHQQKM26tcz2Jcb2cRQiFQdlGQGeiB/3jysjcg5VsHGFA1xzhQZt5o3ZdPGLpi
LqZaQFGiTVh5Y96dhG845rw96Flf7UIopntzSbpiw8KUKoXWhROe0Ax1FGG2kR9GVIlXJQ8DXjWH
eInaXJHeC/ypFp/mHNwiRHRCzddpbv/ZwJTNOfyzofhfYuo15+r7dmyHZBrgtr0DT7mYQBc0dLDw
ry3/bJ+KOzxtXKO9pXMLBnYKhx3X/BFSv5/9UanNtkb3mfdZ4YT7RghTqq0PDMfApU622mPyMzo7
d5CzD0XNnXV1P5dka3OiSpU/XCMDAeqt+xFUBhO/NXdd2YCnMQ0BvYjjiMmA/L8mcvojs1df19aD
Xz3KoePN3nG116kjB9lFPB7AVNpjCNFwxwTPlT1g08TFCjQ+CWEg2tjqDfNoa8ZtVCY1mavAttpz
ImJ0WFL/RTqJ/2NzdqPfdTbPWwugZrQknBZKvl12EBA7rOjS5k7Q/6WmgC7t/7XcczQJWjHV7ATD
wMVUXlWUZ4k+oqWDaIPlCQHSn9o7nQ2SUqKrUnzH4yhQoIvJzdoRcanUd22QcuOGg0HEnqiHPhG6
cdR2DAQprYfeMlZt7gZ6hISfsa54MeT8ym6XOPeqJ9ryRp2N8oqlv1cCLMD3M8cflpnwy4wIjL0+
iBVCW43G+KtwXzuW3K3pLOiZR7gmbtX8RzX7DCjy9fnHBaUxgnlSXH8J0bOQc8awk7eSAG9KU0/b
D6+SkGTQQQi3cdwfxHPToYkiAm78YIwQC3OfLJ4AQBlYlrbcqAmqdUqteYn6WkZLA3N1pAfOKTSH
w5czvws/fd25uc2ekRlKasNEun1DBSkC26/Df3vKGxE9/yRIfeeMNKcDxmHa13ZoOitHgSEqrm+6
di3ekJlf+kNXTRh4sBr/EsNQ6Af+OW9uqtk2i2Yr0U4209b6Fd/jbWr+pE73DGCeI8WZcffqFpyT
6Z+FJEKGmfxpr/7yghdJNsvq11aLK0AGqodS6iH+FVOU+Oou+bk5SfaS1hW9A3RX/b/beLTbI+GI
/iDqZoVsxj7GsFIA8reqLQMEeKYqHqANZxkWATAiFVnxwk75zTrQL+cTyb9J6iKA88oOD8p/8Sig
AmZZX8Jjszn7Dg6nsUJ5CHrP4NGlptx2MSpd/ExK2qN43ZXE9kYJAtp/2YVTbKqk1GacQuAeh98X
NbbrqdlNcoPxgFGYKW7Fan0iodyI6Ts0DjCYDPo25Y2TUvL5pJN6Pl88ezqbnnDA0G9GfWfQ86kJ
L2Y89alriQlEBTDt9VplrYCHTA/YeTXyy5DkgHzJx6IQMSLoLACjPhiicY7UMqGJ/4l4e7b57fPQ
rLohCHI8UJnfu+E6cpwMbziqDx+pxHG956XOH8gkl1/kvRf3SYvlApSJFfUNnBLIypR0qZmIkHYY
hgsHLrUT/Rh666ss0FK79brQ5izh6YwckwTIzsyPtBPjWdwQA4GfkMIEi5s8+6VS5KImF1RKAzQi
j/Olf5HUGWq5idY1aqGKB5yjmafU7tjm/x2BPiMLUK+GYBRTahVFj+HBB7cz/NVt80hz1Iglfi95
Xl7GXbe9j4A/OoY8rGxlAY6Y8g6P3OM+5swBxql1HLkL37BdjswfsWq/CJl4y1GKpTPAvsO8sai/
1lg7Hko1rYfH6zDPYjHPP3bXEzVUOrp3dPluKPw4yK2uVxCoQeeEUSTg+mcFjW8lvzNGKHi20P4C
Vwn5lZbIxM4n3Ma9skmqdSCH5uShrgR9oBxQ0hm1XCBzOrqVi+uXWTxlU49MvZfSWs++mqzwIe26
9Ara7YxJ4dO18Lk+d6ljlli5V1i51aA5Ox1OH6lCreA90AVS5drE5ojIQbBb4ctrqDPTIwq5hOhd
fchWbyC0ckQ0eUyvd8yO9uNs/VeIGFY5b2cU3L6bWxroZVdv7b4qT+TG/AlBou5qTIBXMOgymMtd
Mb3TYBagF6yD3lLkHPdg5ClRsEq0y0JNCFms0BEqN5oaAFPhi5f/N36qwxU7t5rJnGMjKY8DXKpp
LsAdpTvPOPk3H2u97MHEJYZjW79/gwz4vvoqjGVu2l/4RgFTIEHIBtMQtvDMwFvImrXg2rQapNtj
vLd2FBdtLkwrVZLnjIXATPP14tZ0SR8gJiLB/AFcmUmV8KGer9RV2UGAZJY6ROonmfmMzxqPc9fG
dsVa7sTDg+Fr1roxAxhyjy1WU7KItSh77UVkF29rJGtRvERZgC+/DUSHTT5tvSn4xiOyujSNJl1c
1cfj3wgSSfIvYpy41qdw+HHbh1K6EVerVjGyRyxMRHVsLwmHoh+z3RTuRcWTexj3+K/Mhks+mj14
uCAnkpVDudydkbQJFPrlXFO/GkQf6g8yOPVBUFNLVoaJGOfVggfEG+QZq2tzWKjv4uxhlSdNwIl3
rBm3ow6CAVnTYlZlQH/13KSF0ALCfAvRP4IYskZw1RiSH6Xd5/YRkUmENywwl7g0AXQ75fxS1tUa
pTOON9RBxSSYwSlfcszYwcO/+dBF0SI9XoGdENKca7Dqg09OCD88X0vhZNsOUv4nbxs8OjyBiz/3
N6cpHnGcsGsEtKJDovYh0etXK/8vKO0HICTlaPWNp2Gn/cwBPuNDiGc3Dku5DNAhwCtrz2s8rYJ7
+NDwi4SIohKpmUtjE7Ih1qfl3h9A2iQ/64OW6dRgstf03M168y5iGSX5/kXKtkMJXbQjqd7glbZw
HF5JJZtaj2sQnyXV/wrp/rvDy284iRY/0amYawZlHUmdALjhrxy6B0CFDFMmGsKYskg7t/nu5fgG
pzm/1gAVjX7chQiY5w3Sa7PzZ2bjXR4OPbx6npagv0qQIRVFZrs29RJ6FNbnEwtcIPJtW8vBIdSF
gijo3g2kyxepYVzVMXhvxU8CXmBKpBf/9IvZ5x5agDThZJHWx6hXVPieTq7zOyCPYsp9ZDTn3g6q
W9x2AS+y59Mz9Gr9PhIuTZTGP/6rq6mh+PQ5h4bIoELOeGKrC56B2jfhmtufb8rYMActHGO5z9tW
wvAjtiMEAP00B+Iw/m2aT34EFdu/9s1QTCIwj31Eve6jGjDXeJbuIHBa0kDTY8HFfRfT/MXn0vGT
OwIG9d3oJ1NaUT6lIEBNgGOroMcejTKy8Yc4b48MWllrhqs4YxzHA3GlrPWjK9CFL3mJMBH4k6JT
eMzNmJS1XR2897vWcY2A6vyVXYGVz2Se9O/k1CuIPDDDyHc5EmsvqUIoZoXM1/0pvThQwoRIT6cp
pfFt0GKSIVbW+pE8kuKSq9DTqLzeeJRML6nAvEoTKxhCj8fw+Kuq7vctgGPmmu4ugQSteYVjZmOC
Hd3GRXiL2etAaU2tA0Oq8ew6qNfGlLWPMxEuDTJoYwVTzEUHvOjxkDSbtftd8BETnnYgiNqaPeID
i1j13NDMz7Pxp/NsgkgOl8jKdcO3MAaeS8loYV7nOsqosF2S76eznfjr67ueSBeupLV3EQ1lBZaQ
EfzcihkkBHXF1d+34lMoRIqDW2bdNKZQ39TY4PXRYWPseKObt6FGQbBbe8BwtLwfqzHKpC4VEIGC
zkAHizxPoaOkzEILBuwl8tQMGo/aU5r+au99gqzwE7TdTUkerBQ5DD9cXuA2d68lZI481u1POzFP
YfoZcYWcznJlVuXB235YxC4YiYWj3qUQhRak1crlQtDyh8b6TYRybWsLHWDceT4I25L7curKopSS
6QcRbK8q2YxoD0eg9TEW092Iwxn4YLAdpmaIHgo+YlqHkJ+6KegGgoLNdJceNIlNXJckGxoeuqOU
QtbsyqkuUHWyltnKyri6BUa2AedZndhsLe2kkL18QtwTdLUwx+3ZWtJES2ONvsB6FPsZ4XgP9XWG
fYGqASfuQMPySvcEp5F9CvTrf7rrQ4Mbx0FetkRjHA4zNfL53EQSXEEZr0ynJ2HQ+8FoMFF6Ovj4
sQjscWa0jr2VLw2VF4uSIofRlDgpuhxl/oiVdX7UNXflUv1bLNdJmrC9R2hYZF/keRGrzNfMNKft
VldzArgnpI374CH/DMIv6qFCSyTUtAxuz8U4+5El1Mhb2ze1GM8NUbRvb+mQ9mwgx+l2ZX5Pnsg5
R7FcBOTQMRNiGFfPagqrMZwzWhGinOYXxsd8oeR4rQZDQu8jZgRpY3cx8ACw4pkoGe+juDt0qqI0
7UdCJDZ1BXIho3XMoU4hvPxZNxszo6H8JOd1yl9LltRPqao6LK34M6by9D2oVI4Jh5vLCvYGFxY4
5lPF6vXAKRn4o6WrFsL5LFOB9h3vkMOaBze4IPS4CcJDQNWJA0swllQWsfjDTHOdFQswh1DwKh2T
m2+LRrXNcMSsNAtkk60RdThUz71CXuKdJ0i23cwEGuzRy+UU99tjU4evtbIBobpuxW6ygElCHfHK
m20ORRFs8zWtCu8GntOM1NobUc1V/onsWyo7Lk/mCanipbcYzP7Gg8HugOhxrz0rRzXyCq+UBvae
YROrdLwfjMHADptTcDAfA6GMOfWxbhMX6gzexKC356it8YaIVQg8TyBO5q+dSfv/0ZXsZHoSpIll
da4TG1I9o62J3znEn8EwSdKammcAGY/dfU8dtZuvRlgIXxKiFNoDu1EUYYKCSfiVuXCxSuXOF2Uu
LGDwc9fW0Vl7AZKP8pINDV5QwDO5w2p5ixh8r7/7ENHRbXuv6iTavhMKZ10fyGEBigZC9fuVj6o1
hmISQQuJcGNKuAioMgA24MS3HD4X5j00LTT2ylhnq+PRP5xwGWQ31+j201AHS8LUZ4+xaRGkgtoh
4eIzYetu2bkaafVJPWZWS/r5ndDphLEQtxGag9XPeyhIFu3UI796I8qVrkLY76L7U9h6gBcXAFDc
5HVdTcZiAKDpVCl1h9Q0LVYE8SwucckprU/CDuP0pKhTipn1hjGOeXHJKAp1i7DNEHO8OIB7KfU8
tHO5a3l9pVOwwuL5VA7sPyfJGe1GuIrjkGrK+1Rcp7kI2KCX5CgTp2mis9ahZsYBw5BSlY7ldkb2
eWuCEqJAoUG3ATgUjEgIzQ+QWUZs8ml8vsk7JZY5yA+uCeDIH5rz7OHN3rKurFZlzF61GH4FXmmT
5Hyr4UVwCIZOsB5D3Y+b3jlLKX0UgECLU/d+D+atNm4iSGg9PRj2hQbBno9qP2nbqjSH1vWbZk7Y
emXyHkuw6z122L73lzt/zz4msudrOkfJu0uLlAUCqBnWLfgMaSNYeqkrYHYpTY9JvLYmzdJsePwu
S/t32CsCPxUmnW6a3tpzKsUb2pIpZJIkIwVwSuK/9ziZ6ZtrmPj2cMevr1+n3XZC8XLxnbflpOkD
C+ORBYmm6B3EAusFzTSACxZtXQfn/u8/RjxIYmcXALzCAlrZWFTOmK7HILM/YBOTqfDgAq5G2skD
2Ro+ZIUfKk6VQGTCC/gX0N17F0F3yDclHo1PmVejLBqpB0oF4/IklCJ6OtimYpVXsyQqE6ZNhsU0
Rdk0d9gi3HaEjuD3VPv0gosbSme9ug383v2hNDNnKK1mAXuNgALnL9n4ua5nZUIgJcm/oRX5ejK6
0q10c/iqIZYJSl0OQAdxykdZP9UuhS86hlGlcwuHSITsWSlFCpT/Didmii2fu9l0nPwPm49ab5vG
ocqNErEJLWGmvNudcgK8I6tl6/KGiIyuDCSqEjHWvsl9X7zeBxEVGElctiCrwM/6LfWHLOVB9iII
hqjJsDOFOKB9BOkEX5+7jMqTuJa+BkSusxrjGrLjfbAemgywJXNpEuDsk58APu/rrL9AaGsgAAcf
Q6YwTDkdIgVLvN9scmZyePifnA2dUrWG2bGA0jD0nhwCP/aKV85klQjNiyyfKt4OaTZ4qEs6mSa8
7fGfdbjrgz3n1SR2LHh4s6TsDX9kmkIZDmpHpN/ZAFtB0sHcv0+y/7NBYqhEKaM9K2XMnpSbhrt1
jMqcQc9VaTCDbrMIGY6C4kQMWFwSqfEFAerMfmHk+vw0nnKuduz035x9B3p1tzELH30vdyu4GxqF
T/UbPqT8gcviHE7gU/MnYI79HQ7Ew2civre/+19qpHgw0RJQ3pDl75gNk7L8fyazoR5cYnWjrFAE
f0voVDovgLqYjGPr7qTZWpVk2LIzJ+KT9MUHAU1lpi9Jsew/8kDTcrzF8S9sdnRze0A0ssiAvyR5
xqLk5mC1byzT15dUA57bEnZPoUBh4a6Zv3Pp9rVy5h3ZijahFtqk0NJoFM9GmR8EE8oQHCwGNoX5
Cqtmno1yqiNRa5LZW31c6qcFalB57CeQGb3dWrUGMjwfB+ozoNaz5Pw1qmff7FiSNhhDghIHa1eo
eh40zr/j0uAGnqivFCV7iDdTD/PD6XRFXfIhDfcg+m3sr8lzHNZeDEMYlsK9J25zoMMLyE2cZItv
yb19qQ6dvSzxhFrWrrUSQtSNqSgHF2wcrhBWMHA07LRUsTAezcrDZn3MWcecP6NsSEIuWaxmNcOB
ZfX9tvxRQehY+C5dSYGDR7gzrEH3eT87UTu/8SYujQoFM4jNnEtPJboATKG5d3HkQNhmc+5qU6kW
R7sNrs4dKK7outrOWm8VXqy1ZG4KxzCaUFGksag95L1eHOxGHrtN11ly4uG3Hmmb1asazi4r7n29
ITiDAa0sgP95WkjCB40QWjiXYMnrg0aTdeVXvba1nRZOvlfsNY3qXrzM/hhc+wp38PrvFR8OCO5d
Fo37hAYdoxTVfyAgsmoOFjn6C6xshZtPnKRPRJKQb/x3aXqKSm/2kzr14Ud4it0w0ZgeVMW+Xynf
aaNP7MUhLmzPqYBf6r4ey/ILaIrHdPTqApq7P8NOUD1avyZ9rA3BHFV4SN7A+T6ENn7br5E4oJwy
lFnu2lcvj0gOC/blhhlyAxtwH/CsvMe/Hez51DNXe9gfbKvC9ELeoQkCO4O8B+4xrBMTXMdfMm+I
BKijeWBrRRo14bpcHCkeaFTzGgVQw6T7lehfACIsH4Q1U/xsMnmeAwDbaBG6HMn+o7d0PlglVIIm
aRgBKXlpLImiTy7pdTSZGBRNCowdLsFF9N8cX9VEX446HOJ7Br5eXZMHF7JG+gecCRxyzfc0lQFg
KLYuTzh1rqm2efT8NQURF0+YVmTbqBEQF3HTa9laeHs7czxQMPmHhbr/+cxGEo/gIud8HOJmICdU
bYX/wkXAqSA3HBoz/PE/GIX9DDvg006X/PQYC9bof8eMsn/0s9/QhNFs8iFKUeuzqYFMWCZJt91x
xJgb6eeIwH9PJEHU/95kTIdWhLPJsgFc+fMM/CLrRwq3ZgWiT1qjaoCVP2YYBl2vY47/fK/ASLoS
PTpKfCNwK09QNvMzYWf4+HwPqtcJ1KwAegL9dkXXAp1nvVz01w0aoLI7FmaNdBww0pdvMZXPq3Sq
+erhQCyhE2dUZglER0jyg261+mF89gop/4QbJHMZY5MYzP5ieZ6Z0dd6Qt8iHvnk4LEOp1kfhXjv
htP5Miw4ypS3ahA7iLeAMUuYCHnsaQGDVkaHTnDMWg8wkLlNMbo59Wo/RR3lJrH7EaxDsS9KJkb/
4uNJD4rfxAIU2M0n8Hh9Tn8M97ULeu8IC66AIjCdulOd2MGLte3maAjOE3BKvCjtuVsaK0x1bTt6
OTxwD1PJMWWGptqEgYnjlR0Su8VBdsxITbpWwiDAVLB5XU5Xiw4MpZCFU05S9Yl1goLLt08FGsOK
eKByfLd9v1reJScznmsBe9wtiqzQLdRA7FGbgVh1UI3SXgxCpaMT1U2yAY+Hj6/WAGVHwOOojeWF
EkS7D3roJL2UIZOiv9mHuHzEI/FEXWQbAxFuyP0+3o3BpK4DlIJhCPI8vevKUIy2BmNI0LPzdnzV
ZoF86KusZZDbQazfyuV2kdSRdyg1fsl7dGUVwUojQ47/pjbkaNPTGusKqzCviejqwl9rLmwjwKHu
8Y7XuSu3ElpN2YeJZHoR28d+MEXpZz1fO9Bgc/QCrnSiC6AgBszziLs3IynyDP0Tzpb6RyyP0hM9
o1yh8qhqh112oPQZCUBHVSyiHmJwP71GkbjJcQYVr15xq0XrrTPd+nKW7P+/UcV3zxi7h7Hke4B4
a/h+YtSYMlpdT7UVrIGLuMdv3QCeJ9Z5SQhQnftGXDbPcIMAYH80PylUn+C4DDum8Jr5pSr7imBw
ohXyB2Zim4FitG8nv3ll65j/PwLaUbla/ZI9doshhVxjmXS4BuTtdP8DGkKUHNi45l5U4VJ9mgAS
Zig/X2eFNHKNXH1k5wISbBBNa9i4s8x7YRBuF4ImoD5n2VjB2ea6kmqV4se9uZ2wQKMsNzeMAzMK
4J/bxhMwaBqITN2Wl/z0P1M7Oa44cXhEziMlytzYLUe2VrltetIGYxkJcyYdY+LvIeIrWXaYvPoZ
TG516wTYA70YmOITbgwMleU5uDVwQySM3E5AXwH3ommbP7RHR3zPtqXk86e5Aie2aYt/XoGTjY+q
dfFROJq4iTq8Dv1+Wxen3SSuCXJHGA1hfq5pf1ToJktbliC21cvpjPjYXBKgA4O54SsXVm8Z47B4
z5jChawrXd92p9I6/ZEJSwLFSPrWcaPw/BNAIAAHOrUpcVj8cK31wBd+WxEdQCYAbJOWAenBNjOz
N3BjcUE8vtUa1Oq9S1h6OTZUwVG4r4Ms8sZvgC0PkuxhTiEfoRaH4Q/FbJHA3EI3nSYNKkImJ4U/
69uZg9lM8zuVLcWKnA0xMeILCWoYeuNas1Or8v07LDoRT0+ntLGwUi57nbWBFG9Sj7ikLhB8zRKf
VpYmTiLcq4aHbttNHs79avii7tMucVNZ9a5l65lF/tYrUmKXDjqzX7ubOocLEUimWTauVPkc6E4b
JH89cnV8iK7LZ9IvXWvr//veBjwKgNwx/lr5ryfeE973jJTCjvbybNn3r6s3qKA1WI7ajg5FPzPY
Qj3BqCZ0/ZAAVF0wZ9DYnJAEQzA2oXlcSoxJebqWUrKM0q0HL2mydeyMTGhZxip49+FAhD3xqfsg
L7Wa/TPdWmZ0gyZec+UikA6SGcycoaAiiH/5PjSEpaEQTHWxPiSe0PvrSZpr3PKU/KlogerRCKIR
T6GgF/BzYYTJW1FWs1Nbi+riSxdSEsfYbtmybozri9891vXZzHmcw5cZqlg90IofFpYHMFebUSUg
fBbS7LSXQ2ssN8ViV8oqkdvmLHxkw1fI/j2/wxhz/umidFubVDeD3FdFDh9NKIO8lJtuyPiMjKQ4
fyFKNDd8J/iIlfg5/O9AET8PSPKW+LKLTr0QfO90qs0minQmffThKsz7UpaN/QWqxpfJ/K4o4wok
T2I587qUbX4jxVrpxKkt3zJqJnaLQ/ergwYJjWQI0kLQwGcPyoggESEmUvt6WIcEDm6GFgo6+SSg
Nr90jmjq7j8bwVZNHts9OTbaQdW36act7hFTqnrbK2UZVQ+edZdgN5vfZv8G4MRXRTDm1ntFnc/G
K7BQ9xy1JWJyRC9M7T+QMBJkmmxncT1biYJPMVXHfGN+3ThYrjwbOlKeR4yn1tjRdLsEIjIhpVVR
zqPo6ovEzbg5ThaORWZZ17hKflLtWzj7gHfCSrgMmdiVxVzNkTn73Xg8iCF8v2eWy3ux6JRDm2AJ
2Kmkv7cy1wgxQdvdhtd71hDVAW1iVrluScTODDNgyqpB3JehB6GxdpZOVX2HYSn4KgYR4/Y76kQG
Uo5ZrHJY/t+Dx/+cKIf6vUb8N4QjnlpOe6diNn0dJliuhA/ETt4l5i7MPAw4jJQcR6EpOnLjN74/
xGBYdB0QdW9gGwHPmgJnVFRCASpZYva4ExrLunNqB9SKZGG2/Qx8bdSDm40H/JXJKIWxloFNcte2
J+f1YUn3M12Fhwtt+YYmZULqJj5y/IJ7m6fvdo3Wc6H6q4Y25ZT3TFPGcNIXOmBopR9etNciyLE4
tVzCtM5TP2O9VzV3ccU1ytelxNMsOoErURfV3tfcZgqDlpRTJ11MOriltnLY7mqgx3IO2fkFl6p1
JPL4xKQ0THusMxjgItFvZvmjh3+68VboZnkWe9+XD4OE6DOnAT9BbQZCSr4tRdH0QiLjPaC6cl+/
3jD/WCZ1Lk+VP3lZIp9FYoMoZsgYXWMgKYAcHIy55PseSaYUTqfVkysD/0Q78cvveUNfc3gaI9O5
gwH3Xe34DElkSMXAVt3M+WWt+Vk3wA0xG+YZtiS8Vee/QVi6mFWu187dN/owNa5f1jNE2aiF+SDp
juyNvERb/I6cveq8VHr3q9Pd38LqyGPdoDY0HLY8nORKR7FckL65a+5BwOYpkhEm3gUAGs1hx7L0
9YIB9ZizV97WJqoZLmmJOhwKw9IbFofN4aD0zDyALotT3Fm2ERapyEpsFin+SHaw2RJ/FybMvMX0
Ybcg5v6Xo8JHe/hqA+ZgwKEIGlNZ/AQdYsixcaLJOZf7UwtUrW+rWgL3eFd913KPmrc1gIopUElH
JjiJqdKlcUk6AqBYl8lCmcI+jF8Nl56h/U4SAk45yLZH0/M3KbvlsJvlexaX0aVGC4awWsPErbfA
2eTPcbAGAvCRXFQ7Lhwl73sfwmwCP+yhC0FoPKVMORIS6PNkAXYMMbk/QYxbiUct+8Noe2yCk2fX
furzfuIpQUny4xvgL7beMf9HVVMm8tdnq53BCHUGtYmsW7/Ng3OP1Ii6PQP4RAOqnI0tS5G0bBK0
SSq+UEGPd5WTZlcUj3IfPxx5+pL3yOWEirPoowpDbkbK6u3+FqgYYsfH41+NJfiei7z1P24vDbSf
acDaTrEPTBi9K8s3XsMIh2fO+45Ffe1Z9INlEjcXJY6IZK5B1455kwi6MXO+EuKvUWyySiuSk+Em
1yFTnZxiKnppsGWeloGFBoRDgSsTEO2xN0xXwRdAfUQTPsGDYE/NupK9ho+G/7OUO2SrWkClW4mS
70jDyleS4FrDu0XMjnEDgvjqgN+RQycMtpgMRSWWOIRzEMFVm23wqbW5FgaShkYOOeOgpPWUSmyZ
RofOSLQeOvT7Hb5nF+uhR+3Z7Jjh71e9ruAdjB0aKmUmPP5QF1L/eV+iX7Z6iI5bjnmAi7Yf5/8/
k247bZ+v5TEjeoYWmJkTQVdKEQMyidGvS/d0YG1K6trsCdZ5eaGfXXTPzOvKUA3D9oSaAKYEJ1xo
k23zOwhEUJsV0q430IYGTp9PiwBmqlu2yoWx7rSMnTwjwp0Rs4K8bNoq3uZBHOauyFLjV65yob5y
yCT8CF3hYOk2QQgp3Zez/0m7ZMDH5FPJ4bIE3oG6eOWOp+1TGLxIp4+mrjeV/kgyw9a3jB2qvUNK
D34mFdUFgg8TWvn8O9B7O3vbtPv2HITdMv6EReUHPdD1SXPL53SepbKe1JtDQTqdEhMGQq5eIgH+
ipnepfXbUYHRtLqKlPF+7qRLlFrvE+5EOfaYv6kgCnHapqfWlOOFD0YUvuKeEqrAtsa/lE3VemRk
3ga8ShlorcLTBr2n0lCX1D03tXftPrEZZCyqsxcwNpLI9WY5xTkclDNilvp3ejpP0KCTFFds2P/b
Nfes/d5bHDhXl1HJbyT3RyZOPSPaeB1eKDc7MCVojVHz3qDJ3Yb4fnDMMuONgzcHktfQZAD03L5X
z5FhiVHUGBVCO3qfnFgDCWD0Bsvz2/B2qdzvSfNaHBltv9m+v3Cwdn10Rgb6ZskP7B0WP4o69kYv
eRgEdPue3xNCUIfiCxydeibL/2pu5SkMHACRmXmhAY8qwucM9PXGZnu98HMeLkzdMos07zsCDkHe
EE52CX5F/PZw1PwQetIXlp+W4fJa43hORvGJFWDvgpARoU5Wc2AK42xZh//IH5NYo5/wexlU/E0H
K+N2xO9kQap1UP/7jXTJg4Ic1yEPuzR9Sq4zOqduSxsja6PYtWQBZUa7gdjfhC5MHB3nYWI4jOj0
6A30wCtruJJ2XY2Q7xc3MImS7Gk7WQM4pJBLH9NHY/DldEvLxUge/t7hOt+yBFlEocD/H2J6n7DT
/Q+5SzZwix74uTmpJww2uufEDK+SQmMxSG3w2AqgtLSdlBa1xq8ZvEclGpozol7NQnrb08fnvPh1
VcKgynB4HWZTIdRZeRkOpWmzbPzKOXsGedZ4gk0vQWvshTkkbKYUcEEgTleOUJbkMs5PVuyEesM9
Rd6vm4FEh30+dDoISOAhunHB4NzJLt8hiD61lV6HAelxXZrcaaeujODJuZtJGDZuGB/rHGIcl2Lg
uKsCYkyHAOkdLjO4j3zZTn+f7gs+UyRNVyIQe02nI8L2nBgM2HGeK8+4HUUELb8gky0hyR7u9e/Y
9hYw7a008IbzmejywqYVWUVdZDhmtWwsMVeSRCc/dOpgp+pN/r5/IXKAizrDJqDrqnSjZDFZWYXj
rAOWmQLZDBknJ5/Wp1Z9s/+LBfxT538d9WGj/agz2jixszX+3UriwCo1alkU/LwxPu2KSWf/cF/n
r1BGgFLd/Nu6LghLGaCr1ihBj7+418xsaz32t5W18DbWrWneUeyzCF6GZM3kpUjFq/PzNJ86Cf0L
7VZM6E+ITUvC1xAGySzVGyD3WWwQ+KJgcRkLhoTEpHXgI2EyPsvNR2g95dc1DAlZJbTmkUljmcct
/6L0zdlNVmXR6u1Z1RVIz246nd6yWd5NSispT5kF4w1TfUBhRHHFEcZlV09Avs0kzcVC/Onfcloz
+to85AvgQiZ4iEI3rShANfYd6GNktxL4iKRNT5GLQP8+2mfV0ft7sx6FcDDujvmuJ8Jshv+v1E0z
I+xBq7H26CrJpZwU6RdLAKP+D9WQuGO9g2/EgJMB/YbvyUzrqhQ+14yAnjbiOsf7Fenw8m+Yj/AV
3RSloOCBFd35Vp5Ey7QkYVIiiGW7Vgvcwv1XGBkCSluA/OdQxTK7PBZuA6KHqLUXxx3LSPYK01vu
s7LjqKjCllR+F+kXfBOKNpmwC3SoEJDbqX8grubBc9SdujxEBZAfBcLWZIlCkK8reHjf9H+ffP+N
LAjlNbnNjG6KBuBeeoGJaUs9GvFWrCaTGhiBJDZFuG/DRTi7OQ77uPXUH6mkVNn5EtT9pU/IXR+K
39f25VX5Ykobczrx7iOZ/vS2eEwF/yfjfmt1Kikc/c52XEoNYY6cjVZ3XrQa3ofURLlBYsnK2s8R
mxTpQwsvh1dlrKeJCri6zcNZUZgklPMKKwt9Cf/mGy7LnXGhcghXHR6ywv6XLipdKgXBnjepfL0a
7d59rMYKDwMdXS4Vh+fT6rAcnG5GrLAZwviomNfLVQO3KkdsgWwOcbql01UIlXgaxsnaNq0Wz6MK
AHunz5Pc5ZZ9QuJqh38rSj59gvY9dIGN2H/cE/HP302wyZutj7qPa22AvWmXn0CP6cyxkBtIPNRb
ej7pY2bzUA0K1+CxUkNDcFuHc6kip1sW9EJvaQB66Ya0kqiyYj1lYQxkuVLE075PeYtxQ7VxhMyy
tzWDCKj36+3xOA2asNiAWy/3N8b7e9mHoQeRD9xW4vuEsoFPgRtr34S9fj2ctKotmVzIz0LuqTX3
6a0RKTwKswNQZZ9s5m3H8CdysW27KGpO480btIhTuX2n5qiHuKi2wZBFj4EbOds+Je6iQb6sGE9t
wyNHcq73qlQyjz7BBZZlKzUSR7TZNkeIZ7Q3CGjkPBobalLe2sZHvGwKWbL5w8hZdzsxq/xkF8Kg
kYSAllbWNmZaGCQuqAzwIG6dbGxCKSPT70HjFs+zjbcL3BP3yJa/ETTcGmisMC+Vj5IQfIolWc4Q
mutPV3u/x4/F1/cA6nOK+5CAmx/T6g9MCSX66m9+jrH813IYOkKhSb6afnRqoFPIGyDm66JXSWaV
kNEPGHkEh6+tc/5Yg3SwnC+HjIiwRCm1ePb8h8j1+vNZ5vr8P70eMKRr6iJFaJyCByeVpiGeavMu
d6QfHZ5pWqlFRbVKE/i4XcZlXE0KagGgNl7eAUJaoJjRH6k6RcbByu3uObC04lVV20P+a/krdT8v
CSIsbNGBeL2ma6AbwlwoaVOlV4r9goHmn9mtbjWuDorSHUu1r4XTOreyPHHcmopRNSiBiLGlzqLF
BjmhGrQwie93QYCjIV6U3qLnRDEqp07zMdd9goWGGcC1vpzsPb3py07SzlQjT8CDqX3wuFzxlaRH
KkxiLBa4kEsIJsw/+KhDbQjfnV/IC09y3Nt3rNXGVw2/M8HYtRY0zKV7qKIljKbFzuXNKlqlTqc/
Ev48BvLQXeYoIHJOZcClyl6A9ZmOEbR71gB3+M+nUs4QR8i78MKx0pJ7xbpg3LyJ8bEiZ/Rza8vi
wcFVU6qD30fy/raykCrOUujMnpwGEUgZ41vdqUO00bkA0LytPpgVYFrjCNw2llvl8/T++poi0Yog
SU/DOW+xs4uA/173Ap4Fo7pVhqwape0IkA3wHIglbSTAqwsH0MCV0cUPFBZC/gNdD1JQNU2rDEwm
6RvBrAqbTdhTc+i863mihsdr5yJIt0Yo00oVa6yUAKlaQt6gZaG2fsPduJ2kUwFNnyHScInpywto
1kv+Pozpyme0RFrkzynXtBG9IjuZXGj/Mci9WJUtbEtuXHPQsgTVCmmlhGBZ/Fari7deT2ZR6WhV
3cVwKccylK+fh7NPT/YmZpDhLpxF3IoQDlQydqA7enFRA6v1lunoW5iS4jw2U6fxLhd8X/+Y7/eZ
+gR1UrlZpPqLBkQA3F5b42QYzg/DUCajBUdb/3jBz9ljOU8OaChridGaIdfwLU6yyH44CX10VgBQ
lH4C7Nj6157d/lqwZKetV+5NRf5ehtXuMNnShhR3J24/CTm93PJ2TDOJSKXs7RmjPxlNAI1t6I2D
T0Zj8cwV+zYoggJ+mb3QqoApLp6sMmr1yVElKZqjBfzHOUaEje1sOE5poWBF+P2QarNS6Tgf/eoL
F8ZN8StH/6iwQuHpn4qcHGq37cjFmUOyvIWFiqoRtdKTWn24Uk2WOzPnl4Sgp4vR5ntfDoKufBB9
w9hsUzUbc4jzSiqkCULYugagDZP1n+fUaeWRTTILWft+bKWguTgnp/cKkfSms/Z6QKqEFTs/ETQK
ZiJlsLo5LhLcjCrjfAl+V7cEdaek8xWufhEL/giH5PVQFj18iI+A5RkHFaDlqFHOl1dNa8BsvXgZ
Gz//gvGcesyqyhFiZqWze/uvk4hN5QYqb13CDeoa9ythWDK1hY36pSd3VlNd+xyLAi+KPQJPnOML
/mMqyGUefWZ+kjL6WqNtWkvSGg4BObKiNFUzT1zDXbSo5reWLrOc/6d5IsC2gFYg1G5wS/I7tceW
95oksBgMmk0/ycZ05oaEDEhFRR71aUT1kMlmuI/7atlZ1cPbD66YWggZeZkJN7/rh89ueT+X3U1q
8ICyQDObcaSHtQF4GHLZpq2UMlmkhcm2DY+tqK6WGqbI8Hnito/xZF1f/Es35KNo2JLggtbeGJDq
hFV0GHCfxCSxZ7bc0Gr3nqxohqH2iNj+55r8fwP1j/wWDtcfZ5NJHKDvhsBmTyjL1wUgY2PON11s
8x8kNt8zfq/KvQ2DnOgyRpeN0CcPsoHdO4V1AcXaPfvFYZhw4aQ+PdEnFuw7Oujg7BuHVLtW9oxv
1e1UFpsUA1XHum03zG1P5Gbi29jBmNG1HbFudBQKe7g5OQX8rxFWu4QTWLsv7XDFBVeDS+uD38Ly
bjnMXLOvyC44N2P7fB2u4u2adhB75pPq0CRt+lr5pRHY57hGdcrJjWutx6akvq0SxnRa2jz0x6wt
NQAHSLOZ2olP9XG8gcXnhW6qjf2+LMFe1DNyIepA/G6o9BhEvERsxhO3Frf9oddMQ001KcEpaKMl
0nwNCOdokWXJbLU1MB8sRLbNnusEwIScpNwsHoE6zlj5A/bvSBG9kxDGYAvc3wLexf6ZcFVPqY0D
N7YUXMEWWurJS/EzBRg6oq5qy2R298cO8HbpYS30IFMtLjAvEefvvqYBAqzALEtOmp82ws4SI6mh
1Gj7iZ+ktJnTih7ol+RPuvrhYAjXCDcjISM9hER0ia/bXh7qWbbs3SHFffjMLL8PEKRjYYMwhBgP
jg6xZfky3QU5ql3l6NCmCEozDWAmtlFgRPw7iPHy2qhZoLNspD6S86cJu98H8ZR0oDMK+v/q7OEW
RClJr5AXu+fgzmw3qxY1FJy1cAXy/3bx+eKmN7oUkCcf7YR7+iuBXHf+XNyMuK6BMKNXOH5BjytI
P79XXqw6oj4M79eM9QLNK9O/g3IPSxhLyX0ENO69bA/dSPrC8b5uPyBhsR/ndmKI1hje2meaz/Xy
czxsrDgqHeOMzdjeHxymqIhf23mhiuggx1Tmi6xptOLWp6rwt74UsQjT6PlZxFPaVIdtYAHnL9yh
kq0UQb57TlcTu9n9dftI1DKD5eNJ7iYZFXtt7ZcCI2V2Kpnu/LqGIFN+niJO1UekeQTuT3MzkQiE
kBT3Zmz2JbHw00+cyfuVR2hx3pjdaZ1AHFHw9lRY5eVvJnkH3bddTdZQ2C8sqAxFeNETmJY4kSd3
PFyVzKpgTJUprP7EBzjPQIRRGQRXGYLXVIhcipfBX37mG0RGNZ4rLiWC3UTSYd58T7TmgckMXZ0I
HU0TjMTCEw2NuC1bLqPQ1KTs9sS3QfAxnVSZxStFB8F9gYJ7rVMnNtG2wCekFiguCkgLrXX23Miv
h3YTgY2vuJAuHbRdW5hgIZNfI9NnR+r/94oD/9XmpSLCmN3X/NyrOiUjsRCxgUceF35E6GGIskiS
LwZJx1KMZpIdhacWM9ybBVfqV4j/riAahuEEhQvkp+U5usV0X8VHJpe8uVnFNNCtG4aDYoEpUg/w
L2Arv3yY2s5vUtrpFLt1gAzD1hIc+WwhIa2UUJrAHocNdDxUqDJp/LcCOwkzirTP2KU4tuphEM7S
TKHgTMJbBmTjZKEyQ1GRkrHxuu2pdSsqlAX91ndXBm2Z1nPZLD+m9yag2hDTnu++yl2dG+YmAkLt
aUTTdmLAxCEj9RwZWGz+qtd1o+/sQH39E/WVKKlbFkczqoCmxJziwA9+JUfn/+wKRQgJRexsw1Rz
e+xWs9OmwTKJ36ZUzKhpDRbm8Ctv8PHHir3fFsW8vkdvYxEUBI0Sfa6+YcDn/SX9aGqfZIi84Xkv
+qbKMS05mp6Bfz22kWy5ReR7r+/sxZBgTrX+cwoN9Zk89vKjkY/lgZHNHYLR4cXzEGYzOvr7VHQn
bYDV8PbjtkScJ7EnsKFwGWGE5A+WAzFiQZweHu6w0XRt5iOSpAlc9lQMmVAoe/BDFWn1nbEPpRfC
lmYyAR4ZlZGOCwwnfrmCGaex9L7WHleE3k9eUADTtlKRfq/OvqmiSmp3+Oio5dbtmb2/5dPT6ZQf
8MOw0ccpp95FMi1J7B/oGtY4XE+Zmk4tZUjbNtxcsZ/2+e8dRwbLzLz9p302mYdtpw3s980EwlGL
BoQCvtgYbUptQTjLjbYTN4VZcuOSgTTRcmE6iBtvc1mtMRG+AWNfYMYjoxcxR1rUPMokERnTOeQQ
60Yx5ZPCz0yyuqdEcVDs7dB9MdUqTuzpMDb+yT+vTHCHsIP0Fud88P4BsDjI/Z2RquBvyrXUyVR6
kpwA3Xyn90ArCoZE9fNgOSCL7KFS1zVJN10UGJXsh18FXdW5hoWanQULSI2FgyqrcpDbbfHnrjlE
NbaDi3UaUSBSUUWI0YNXzzKcZAEdeeGIMVeptfHOjUO8/FOAL9x8hd2XKSRKppYF8faBNmyW6kCk
nlLXqDGB8vWsRaYtkG2JwB4xnaxCSAxE0zivD0EMVQQbdjs49bALLk2jO8ksBdiHvMK6fzANSpkW
D3c+V9kN7lkTXR0uKMZ5v8KYIj7u947NXE48qbCKkQiQX2ojsHFuq2mFnRgov9pkqTo8X01yK2x+
PU/WWk7ChV1/gcBQIq/FdeQWMDIWP7hix31f08vTLMK8anvAMH8EbQO8sneRQJWh9Cj/tehvOjnu
LYcio4/Y1JxVwB3Lcjog3d5dO/Hb4/EJEJ0r0rZB3CYTjI9aNOHVNaVHd24yhMJXFvnoczRbTVkw
niOhdCUrXyBRRuZGL1b86NKpv2beUbXr2LbtSj5Ymo6Xe6Eg8AdufRDkN2Dg205IqcFyz42HQXc7
6SwFapNnF+uaRmz06ontnaHXz1dQu6Tdn+SQIXKK9dYNoEsbp5SDYcwGDtJeyBBKN3k5H/33rOG4
prPiWJp+7vH2Fl2BzOId7qONRjXWi7k0042dnveolO0Tj1bj1JWrEWQfw8KP7lBULsROa2PLfUzN
sngc8XL+rTQmPeoEn+aJ3pP90wJNcIAuUQivg2inOb4kbRAbnjgVMCeNLXrsx6zMnM/05IQ0gV/M
2F6HYwVSbD7b2WI0pMhaJX38fiuRAZL6QSFyVXfiPvOIqUBfpAKHv/kgTEpb7smm+Vm5DYqZgEiq
Bp+3ap1RHaRMe42YFd5BOIKnU4fbvobMY/SSwQZMQEuav4+qSM+lBHYwmynhTMNhaMhae8ejDUVj
qPmEYR4hBmgDOQjx0zHDUQo2lIHHPfHkVoKurs5hDeLgyzh7e3lGvdbckHZwPGM94/84x3RvV7li
jRdZS++yVdvBa3QnSRoc0dy9Ify/N87f0dgUZo4AUs+WD5mgc2QdvgR4/oCydgxOCZUE8M5CFmj9
bCE+0PIBTbsy1go7G1sK45o1fb4YtIbdYvzQWlTlz0TqMv5nde8Z3mRr21UN8tH1b/mV8pVgpqNG
K3vk8zvfcFh7wRkZxr+s1aDceKhKtUXv9G4S/a86csAgLjbAUlLgmcwi1rzBp5/OzDwJBs6sSzTU
tFf3YfONhg2L5EGVI18+IRXWACKaGIZASpDcc/qkGC7slj+c7PjxrLSqxfU3qoNaYhifWSMMtEYQ
sYCozTj5jqwYRPwxETRDU0m8aFENdpfy8JFUjpcppzA3jyAjGLPdzGkQ43TW4dBi3YoAmHDP7ES/
NdHW3XMlfBuoC43gbJPH0dfk7nBfaaFQ57QyI1GaD2tQCTxKZqh17US0m5POeNuTVfr26VuhD5Dd
Fi77Fl6ADG5rLH6JoBT6/8q/4WW8cCIXgZttCgGNGY1cZbsvEyVbFcRg7pwbZqCFm2priVSTnm+s
1TZtYlmhNwAMEO5G94MyB4BnSKZHgPV0hiljdfnCOYpq4m3xwFogLKIy2jZTJ59YFN+C5Z6EwBqw
jZO7MhjpIiYcBcmdrYdmp2vu54I0gaWWTiTg5be6IGVbmbd8iGPzgm5JQ4yExBaROaklVG37MBc5
iGpu+lWh5avtmmarL94Lj1pSY63YiZCalT3xmUwcVrhHbqO55Zt/BzRsbAjf2fOBs8bHERqClEk9
7mXWF7kH/kY7eije94Pb/PPdK/RMvND5+IevMoWc8wJp4ls5pHg5ZeIxvOkHfi+XET9t+BGek2V1
d8Cp94Zc0ETA3pKD2hHpBwgitOSP8K8bRDv/PD9uQudQ9Lwph9eq0e050n8n8XsaMBp5+T3znuSf
GFRVcsb3lGe/19d4KIF7f7YUOPQIXvlk3oIoQ36RBXQLFfLWzaVnyPq4wV9bSEtTpgw/5f5d5JPY
pIIVhatqbN3M20DMuQl7lTOt/4WJBycbqsfkACSBfQy6W+UBd9LELLIZ48K0amqe+ljWRBZDpDCB
Jajh08jLm2OOlGFALMaaZ1nZdsOAFIK4zYmt4kFAYHgHGgA8I6n6vferuNwc41HR196OSaXejHE0
+O4P/pVTM+ycZFIyIIxeoj98THvrVuSmYMyEhpjgfFBOthadvgmHifQ+FobEnopmRV3Di9ssUJFc
0ENoTym7F/k0dZh7qdySzV+lkhyFRrCK3ZqJXtI9guWXrQB8yvW7vLqlcg96QCbnHT08vy4ljTke
TpWmHyNM6cXsKiqUodHTrYf+zraslGuwPKsszq4KyrlJjsUOCuvSsCr2hFsbKusfrwtAgd8t3Uc0
Ua++MigwsAdXFgpe/fPb0EZzuDEm9hyVD6BLY0wGrPPR2EfjrDSGn5T4Ipv7duhVXC83yKWkfk81
p56Cusx0NwDcs81CXunoutOxO3owZ4FCLNFqsqIBNFomWYm4YTsdmy+i2xaHGtOEw6/u0a3r8nTP
xSSvbA5J7flVHJjvp+CwftQTw9oRyk6PyL0eA7K7VO1q5Ug0uoxZo4V2bPt5fjPclyxFY/rUCXoE
k7WqukoX/mQAaoGDw2plG6KGHzy9kyiuIRmBxwIvOREkjx+zZ/ZTKwwvUHM15MQe7+hiFcKB8wn+
3iJQXkCvzPuTxwQWE3IqW26uQFoS81g/hhFENh0x/WqqKdRW2zUq5tCHQeXIo062SHqfG+8B7yMX
oDdsOPmRb0pZdimVtqt5qujWeN+BvBt18OCHTUzOLIb6VP+Itv8jwxObirEs/iEhAgJ/5hi86fuz
BSz8wMiwIIszsS8tpb4jYl50YBgsVGYnM8MjG1CQDcQCUmWMFHOfpauIhA748TRXb2+1q0W03wWw
m/3BMuV41HEhsg5tngr/nPfWuPBE4JV5I1Z07ostZcd+Ni8PABjqK37Fne/sr8/4zywafs5M6IHW
6VnosDyrDmffua5Q3tL7QnGH/cUiuPHl3Vrmv8Nj1jLkqI0hczOPsf0bKGg0ZLkIdeiFFxX+aLXH
T6tEJrHGAbx5OPCQUjO6/SInWqkj5k1jov9eS8/ANcW97eMGthxhQqiHA87yiKhAxPXc0B36RgSc
JSwBds84D8VFd/zVFXyiRx2mtGuunWSq7549L191XQAPCM+D8MHf1sDK6In1PgwMjui2fFhqEONH
YU1a5KjBoNgkFo+1FAww9u/yxZ7pd1qUBOWanF39D/OI+eHihUfsfpg9hEr/EKnKckIKNL5UxBmz
NwUxsW6J71cO3F+M4CwKq+5XNfWFnvaGzGps88NYWn0AQ8d2LTAQQHJimWGOXJiKu65o/3ZX3kuc
HMpuDZjZWAjO3AVr1/eQrDSp3X+0/fzfSxUd9J0IO65zZ34OfK7HiDl2eqWySkxJgjqvmNmjaJvt
SYXqRxa8OzrYldGl37D4ZPJ+5obvfHO7ovte/JsdvTi+X0NTJvQ86LGc5+cbmrNn+TqcxOmQncn/
8qaxDapTH5K5QFWkCaroUWl4GN0gpD3NZZ5PKU/Bb8XdlalupHmDmeFsZwIrL9kcLW2CGQ2itCRS
SnUMoQ3JsH0XZf+5OEi/Opx7VYBgxGQRcY1PWm60UIDfuwmlIwuK+CyoinAWZfnka+5ILzoP1K11
J0R3nXeuQwBONQaRpxLKv6O/Dy0E5uDe6m/5Xo5BiHZolk8ruaBkuQFFKXeoG9ExfEXeSgVe8kCo
D5ZHSYL6E3F8DvZ26bgNJeytduF+SPS5xnYGrEp2c1WLd8vb/MNK3QyPkXIrGfv1rnMGx+rzj4s3
Lhvz9+XHvL6th6C6HCiNIXRBvGz3xG+zFaCUTegY+e0pTHfFTsBHYIW1mzwj6gl0ili3583GJ2AD
f3tjR1BcJTdPqmANXBo0jcS98XnTVGa8+DAXbIeFcCgo9hxbxQod1m9T7d9AV3v+3iwFqao3AnQX
NuBmNCyGFMSeZXG5vlmcahih/uiGfXm4nAizGtaWJY1rPCPYSCcKHsQhjb9Ulf/NhucBC6oZnb/d
a2zJp1gd7d9VCXrUgBMyoYXUbDv8vK9z45kkj6AY4X9s8rl8sLBrmaU17tSpefGSK+Gg97uOmtKS
n/Cuzp4qlgrWxOv7A3lHOGKpMDdJVUDfNxZUIZtvl7VJJCGhYZdn593M4ZxhNEZUzqw70+qyOQwm
v1kXgj1Sr1bzH3nBXfRvlcjeC3ENwm8/6QYumGnTGmncZmpruByZYXqc7tt06JKRAzbRwTFyAlaW
tGX2xDqierTBqFXWO9EcWborSluZxx7X2my5vmn+y3r7zlLp59lBAMAuu/9zoYy36MXnV1tDvldF
E0ASC+w/Vp2p7zUTEgReKKji1Iy1n5WZp5HxkF+Peh5xmo9kZwCNLParFkGdkWtfMC0wl1oQwIFp
k3Afe4XGc/Z793OyO7BLqifi+e4BnapiaFY4BSID+eLNafm7D9ywUvVmhXBHbsPkg2T+Xt8q9niJ
hlJ7Aujrp/LBrT7XGsiTlTbJbj1yZTeU0EU0Utnkdp6kYPmzHLNQKQrjmUewJVJReSLih34keOCe
ZgAlWM1k69/iaIz/X1pUgEplv9JOOw0CIs4K5tSY23HtrpuF928/KSLEeNPP6eOtOA6Q5O/U0QVv
zM5WXBD66traU/QYpgmW/3g/cxddHmzUysiw+lx2b0iiy67PjpOk+IY71w/BNp3L0Pf6vd3ZSXaj
bwEO5zmlXPBmKu2h9Bz4JJ/ZD7aKn3r4pvWBUyIKvib9g9PPR8f5LNDIfydr3XVYjJqvWAlpJ1Tf
wOhIWXnjFH2BTIhLd2nIzvObonFNAjVqNwqNM5ldC5EBdjZlWGlBHUe6Ek6J8uAkigUlZFjZDP3G
ml4NvE0vp+OPxP6Ti+n2kt1BFPYw3AbmH/cvKK4kOQjb6Gct1HOWr+QehITpAOK1zZpGIIV01439
SOXt6IQ7y7L6fIwnGCDsIfgbHNR99VRohxlsdxHbLhJNEqXqPVUcREwzD2nQ/4KlfoRUj6JUbjuY
JQoJc+Nr2mT9lLUnPpUPsVl8bGkqkmWJd2HIFQrVFLKEmkDxX3KhijLPGPLRBvdQXjq2fOZIyrSX
7KtsRMwjcw3MWrboQswofbwQRM3hnY/4H+FKctM0t9xV+8httfrcdOMeGez8ONpWhONKgrionIaM
cDBOFtBiKzPp7bVVhLQ+xEfUlxw3cftJlj5pkbHIVpWYHahmTOOj23BjJndewOQ43B9HaWf4Gn71
qFxnwmTmdH/y2jLP9LY/Lxufxnk4aFujVkY5SPFJx8lYeQuFFQg1bmxSUYuNJjO58F+ZoENYuwJY
t+w2Rk9uwBY8IfmfmyNyGS3eXesGnejsANvJ7eAz/2zkBjG6bzsjcbToqO8FedeINdyPl8RUWFG4
s40OgHiahCFuHJDg36cAfVpZ6WJhNe9u2h1nKojJlh0YXLQyYUA6ZF5JlRavEYkFJ35ncaInY2uC
WUhAO9PmZ0Rx8XySPRPCm3xl74z8+sy17vQ50AfOBhebjH8VuPjzVDSCCT89ZWoc2bVcq8kfdpHM
TeW67VFXgj5qv3t19dc97fcJdL2giiur+svsJwFiuEgg8rU8kkhfWjHs9VGqr8LdJ3K/lvjaEc0r
2L3i5aHPk1YxBhH3iu2/spJUyp6oPCGIbAOhDZ6ly2Cy3aRgR3v9PUCVJk61wRx++v5LtWmEgj8U
LgKZXKvjunlLjlPbDughAQYn6PYk2xQeJaIlHTodqqsjgc+7Rxjeb0D5++FW/zNJVaPeZWzZfn2o
w89C6Jz0sDhb9+DTqEgfmNmFbiPtMmBnMacgJdAGVqXd0n73N55l8fVivwqUfHhXy3c8Zo37/LbJ
7a4RZHCdVjbN+Wlvkzfn3cNRjV4MTYoz/8Z2aWxNzZ+9J4ID1HClopYZeZMZOXCA8Qi66j3nBsbq
STAuvdlsKdGIPVh0LhZQ7L5E64BtZAm++e3rEDCPaHoan6ItEWWbyCR4HTG2IPQG0bvASQcXeJrz
6WBrlENW6pNGnEFBuY0rt3LftBkblDbBJ2ZzXuFJSin7YBzxyvq0lzI4F6ltXeNzrRxl9VocNtQn
e20l7RNBQM4sBvzTkBxKlFCILIrnpoRNsOoEtBflt6IjIM0XokGUlAQnEdIUgrir6RjDohtQlmA+
5kyMXYKZOv0zQRcgGhkprfpr8TkO3BZuE0Xq2vs4zpZIHlHGKCwhEyhUFKnAetmJMlunNJ8P9CeG
pnDjwPmAZTNIo1kLT4h8CSnfW9S9GCYAur87kPZ08WbvrA/taUJ18iAmj9ypdI1HQTVY/PHuha6v
H4/hQ/phnj2Hxf8HImJI6XYoGNqbxNbRsa1BPxXWHwXm5VuzDVn6OJ5L7swZOV0n97WfDNxAr/tq
81za4vXMYVlp4GkWRHlHuz/dOeRilWbjsoaXZwuxhfIeY2gmrVgi1pptQBUgIQtlt/PjpYSLBi1e
bSq+V8lMz4vqyVfTH2pkqS+3Pv7T5cNUMKzjfe3SPcRkkXqWjgv0IZXbbQcX2jsLf5TFrpEUd+CO
q2t5ylamVOrqqhzey76/+Aw59IZvI2cb9P4eIZlVDoRdYkKg9iKEb6e7l3SpX8BEbho1zd1gwiR8
t+3ATKmhjOhtmDWDil/y5EFTLQmuP0HMvOCjCQ8Kj5mb9sn5DmMHZsuTitTWoij499QtqUOrg8hL
zPJTTO/jCslIPKq8lO9IX5KUBNU1jBJ+kzueY+ua/6flP2nFjXiZH1LWxK20/2SlouJlCdCgKwBb
+wcuh/uYQqfgyVaxuf/runvquwzTbDeRdi4ujhyKmS00cUTZ1xR3djDO3yPyVf6msiIQG/qcSunv
gKw6PZ1FiFwJ52IniDb6kxk0UOR3ElysBsGuZgYlsurHpZc1DS/yabpc078/BiZ5RGkQU0i2eK9l
92j9LYz0ZfMjGzLnRTmsKscz91VRApsp1D/pVVDJ/HHZsYgKu1nVTQ4k5gjxfLToM0b1+2tw9lw3
LQlbx9r1SG9JuXRUJntyTr0qxbKLeN8V0bbh/g5VvuKajVjqYJi3lBlWD1zRfhTyBkYTRTovUZkU
6du5rfzgR9FeoOM9bS7Y/gfpzr4PdBra18BZl9i8s7TRxbkRgVlBaAsGYmNJWB3a3yuZEe26fM3M
UBcdvpRZGHOyPACJwfokrau6DdnVG7KHmMLwIRb3NhSPpFgWzoiJ6adUTIaCXG4vkTAweSQjIQ32
whfLQfp1Jc17+vxvvHl58goFFuvidocaQf3vSY0L5/7PvGJfBEdqmM4U0GZZlEoSreL6p11svqwq
4suzaXN7IOA12U9GxiRIytgeCSYxyobC8cPcUz65awRmeBRpIczSoFh0PvmZDpoehzpLIfk3Z0Dv
mhDvcyjhNoyylTTX9T9CrjGUWTSOyk8Nb0CXAsXwalCAaZy95tETZSCeUfVDoCUjwtLxNY+Sjzi0
kVKKat7NGeiiDn+xUNXi580QXw4O7yfJyArgGncTrEWpuofn2aArVanjxKP3O+1P12X3eBOCLx0y
fYeqr3AeyXcP3YuchSu3BAFvnSa8c+k++VnNsEMM4KmMHS6c3EF7guJhq4GbA2ELbpw+VEu+82kr
Chq4AS9Y163YrRu/f1HM24cCk7UCqMNneqzbW1v1ud7Lpnza//oBhkVlJskM00NEr02cVE8u8+ed
I/xMUyqdVEG+XWBDc45ZSE+nbW7fCu5gB8N/HUIHkOPWpjaPJNtpu22ciTybdUssGmbpmNe0ezh5
Tf9/fvDJzFyqlbhDEtldovb3dAS6frn08OI+1jDYnrP73y7HEw7ZA5FDuFbYvTUO1QGb8+5M2HSA
chQ/I+5G/DJ5tJ9/GU/CeWwyx6h/SrJbG2mjr0g+PulOvIu7JTK0nsQPB+D4YnJZXheQIeL/25SK
jQmS2o0wAVbMCxn4Sh56ckL59qg8eA5qk1TyuiLmFGqgFDdIedojD3455IwsPRLJKJoiwHsob0/P
qI9MX+UKuCWHYEaHk4pwTaoxbuAc+LfirePNfIMN8uS3K8wtpQOm4higxSdkYIIAU2H3ON2YF7SR
UQ3fAWWlWEMB6J3lYWhpT2ioWEfkyDjbojIQvBJ1oFa5BWaspOctYWChw0qvE9zN1qtKWr0/E8zD
Y1tmgKdUNuc8jMam2BD6WQMkXyT3hNsi1fV1qVVp8HWj44+oaFIw83v4XdkTrbSLe699i8X517BS
OQGGzIT5DwNiJlh+rk5YZCvQHdg4qflp7lTxrUHrkywyomMIwjolGBB39wlcM9qECc/dCQDgeu3T
QoddIfQNuX3JzCM3eH1nbjP6Q2px6RrqIZmrVchPRgaGi4/4ieagwyM1NjOlTSMs6fQHwuOHVLRF
jhUpVxJxAEq8ECj4wBKru1OS6n0LNSKxh0GUimiAes9vnTJnPtf2gUg5b10TE6VaAHcgvIoo/KlM
U4IoHGWF4fAVHuruwA3u2xBldi74vpWXZW+7S2HHvLLx2kb9gTKzVNR9TPqzNRgPVsF2WCnJb1Qr
nYLCm1tqHJLx0FA5pb3AIq/QheV7Vx8aqSk6GOZxeW3chS5XTxPLEtdZcFHV9vyquQn2dlgYkZyl
fDl05o56rjwF5aVg8Dsq7F+2xASMnmsV+A/lWPqoMkXRqgZBzcYk4yjVatvdcj2GoStoe7gzwPRi
T71YyE+b/s5ZTrbsr8EGWj3gibMqDE4AXGm2zT6Z3TSQpR9eoEj5d/zqsfrzqoUWIdfKmSYBsek0
Bc0rMt0pBOfaRJlohRAEDFaHkyzrns0ATn7QPYWCk/AbiX5iW8QLNNtJfHI8DuJ56qNrVqXAJjL3
42hm9HimJ0fQdtVoCPSVXCPdHwDv6ASlsdpxELiBzKu2twFu5EBLaoIHm6owHywUqXfYszFgvyTp
9YqTT7HktbXHQQJoHmjhGZldjbmGv5Hx/6OIXv+k5EczA78PSvFpXDVQTc67xS+Y2LdBY6GBMMpp
HnJMZizETjt0IG2V7U87IZoLe73nbtHNtwVN/5Y1HMs3RGDthUcwpIOFvSZoBapyHrTfAuskvACh
kJEeo1eCbhHTm7JgjU56Gb30wJz9wMSP8rcfop3wTue5bZEY70Y4Xd5xDNwRoW0VkAPhjR3eAnrd
q+Sd0JB9l/UqurLfHt/2deAWOAH3cHROSgwnOEX1JOtpDYHDcUPM5ieVAmVgHyAcua5X3rpzKAdq
vl07hAa0pRvuvM02+iDKXf86bCebS+KmHjJTczyUXJvxppiFT2auTCxgHDjEgx86UdiFX1qcidTs
Dr5H60WNj9GJmQeQa1ormvdcpidVnhxfZYEkiyqXML2jkx5wdtVz3rHGFcVCUhiwwoIIzKds0N3/
1hWFs4jxrSDlbOCfBQZepeo3tjF9GfZ7VQZDgvdtfBT6Abn4EpfxYj2zXHfhmjU3k4qLWg0zDJHk
4iif5mI5HS6p85AvQcHfbtE9Fj9dSfyo2znof02Mpdfjhg6wkOAZBxjFdg1SLVAx9XFZXOByKQ/H
PQMTHdB5L0IwArA6BHvO22jZpYtNwqGOUZRUVoZFVbZjL1mwx2prMJCMOjr41h36BgHPxiIn7zal
+DWUp4BXduFHKyom7F4Z3xKsNcLi215MF/J7wcQOCj2gTV72/xTryyk78k7uxBoZwwyBscJSgMti
946x++BnIRDQMKmC+pNSDhpz77HMf8tnR8aRNU6lmOZs7+/g8beVAvmt58gus2Bl5o54l1vA/ZHr
q2joTWe8wMxMYfBnIHRx8/rg1MilEgWom6NPtpi5oEaKP3I53B1rZDfyle1SbaPWOw6RASVgQksi
OossS/wke0HDuveHuXZZIgABI6CSptN/XXSSlQDiQvT9Hexkk/Yw1F7YJ56Cymbztl0Yf4VjyfRB
B7pbPimolHSMLKkEgGTCUwknOIW6bZPwx76kpSEFnqBQeLdRCLe6OS30j3QWnUJSX77vzmlDe+QW
pJrQLvw9URj+ZdnEOLGZOcrPmyGM4+4N/FdjjeMsugPO1Bp8i2NlK6B/MlHCNkWfKa9Fx5aR9150
assJ7FU7d2hj6cq7+zBm6CyCy2quETqfc/d6QuWAh9DIIFGLtEyDxWtjIvq7u737A3tydkHFtjKC
BVmPsVkxJfMZ717LjmXbscXBK65RpjfDsQ/FabSyy2eGFA6BFlLwz91ryK1iNTnb37OapWHE4/Y+
8vOCwRQtOZNluAmduPnTTA9OHrFJKvfBo8Hc2NzxUWPYTlY5PDg0aWDxamcHxJdOCbtuj6ejHofE
yDROxxdNTFDbq83xn/Dqb7b5bHsI6JzaRSvE5gmNA9Tp9F02aJ62XsoloBRy71vQVi8BlPjL4o1W
lAidYRnmSgJ4LPKQo7H5OdB/ug+TNn9j64IpbSFSmMXmTyr3al6SPMLpzZhgqToMkJbsK01fmuhk
SvQQw3iYDqJgKLQhs/Gfs8jtAlv80d8Ef/8g09RC8bFpnnYEcLnBCMJkl9VP3I/E7Cn1AIMY3WYH
OVzSRgirDoe/coc1HcmDgf/UStGqbcrVFIuQOT5cTLaNJf1D9Xaa6hucBPrD2VL5Xqt70ij0KcPS
LDRw1P+QRueT6UI7y4BOhb/tynmC/jbf6TC0afzArhPxz5Mh0F1pJYuv5yr6+0D8rNL6sLG2V8vy
PED8pt2MrOeIDlksSZEKz9angzZEsQpDgQ3Ck7LWbzpagRpNIgR3SIeS0jmbJn2wzntbIfCdyA7J
0EqAabaTUYy1RVqnUWSBrZ4a2seOdwYo9jgmvZEhrznmK/VMw57p9PgMiru/7DOrIQRcDYqn8z6u
LQuqNH2WTGu6soabGypz2MOdltndfD4CjeWgIQbJFbrnSvd9cRZSQUsJBFzbzb99M2Tvdit21eDm
B+QHvL/sMFRU4y/LMfutOD4dZS+kXnUVv3jfFLVqDLwGCo1Lsz/udtsVRjkHLVjjiRToic3S1pfu
gq1wmrr/iSFYHuPEBfEt6UbBYK34D6B6FY5IgQ083ZjOGCRNeMWsmQx5NMM8pxKba3ryLz25Yv82
Hr/IRMTBA/J+2Ol2UkUcGStK9PQzhYQeca+DeXiNqe6g88FaZ0XetGSW3TafEP2MWQtlzw8WZnmK
wf9VO+osVXddhxGK2kHDKpeXjqTBkgIySMaV7UvkIw36v9IRSLczebEL7fYqjOxmzE1QJDBQJYsH
kb5aPs/yHsbuhWH+xaDnOvdViRbYPIDqEgNTj1ZGE2QdrtenEdwgFe81dfcjwpx3P0qyxfxAlz9x
Fv+SaHEUQRMR3YPA4/6ES9+wVK+dpxe59l+Abu98YkvoR6bu92kpgKt+jA3MNmAmEMDyeCuCt0Vq
pvMWdfu1lRx36t8WB2NdctGQgi+JQVAL9EqCyXo22cWcKsqxUM7YJ56dlO9zaV3YiJ06ZD8VzoeB
3ENLaFTfSShX8JjrXY+W//AP6/9Wl1BxeHLEUIvCe0p9Eddfw2cRfh1kcCAOnw3OjTS2yZLJzuAI
8Ir5tFpuS2nvlqg38c5UBNG0UkfjovtRKPiabwE5lzyYKBgJ0d5HzTpSZTHHQGdrABhd6JPIylZ1
rrG2J05RKXZMMZHp42sW5fTRMrnco8cogRpNuKCLU40y+owHMRxSQyn+5dqA7t54Yw0qq0lP/UVu
X9Gg0asVRka+4l4DuLjMtFgwIRh8nHEbS6BKbmgyKvgMIVz+cIGm1bRxA5O/3M5FgRD7qK4ldGyb
m5AOHMVFrS17XqtrZAGIlqW/sWGRZNuX00cIeXtqz432qoV/DLl51HikJve+zN5IOt0eFpwus7kh
iLEkp3/ycFLkX9v/gy0kK4U+p3HizpCJWz6ce8spth1D+6/NIM++gqZQQ8O+D+fKg4BK10mHKbvA
jUBSNZZsXZWW6mYCQ+sZLPB0jlgr8x3lVlipcxcdfRbVIXzO+3E3p36guGavAd6i7YxrpG1Rywlz
CG20CJqu/Qdu7bG863BwzeWcWgHr64qkoKWPxgeV4BU5KLI8tS5vOor78G6ac88lAGAVJ2TAN++g
yJJic12qUOxDg4KLmYW2o3ofVTTYSkv9sbNEq7d/hamKocDJcIVL88IpVJlUUeMq9WypWy1VM8um
RwqCwCVfOWfkke/PEm7Q7Kug9iy4dML315Q0F1rDqRb98/tAkzuFkGODyTn1yJtZUEaGwaSR6yjV
L+iqmIMjmh6NvyIy5dkgZ+BpEFx9TcZSUlsfOiC7HqgvxJAH9d9rznsByJmDGUb3kkxpjyAXxIb0
CxPSnZmiZnVEgdsrGlVpGP0VcsP93Xq3nfjnEj/wp6y5DzAqsZdRvC5UBT3/UU7xMzSBKSj/8byL
6uxDBYpx+T+qeyd4Q5JE32oPavUkCNZjd2grIEmiz77bwuve0aVyycOsQVZS/XgT+BQXMdhKMxK8
hsaPwoYpMy/SPSKhl/U9Jazik59SVp/bjnKko+MOx4mFiE8Gpc701hYZCUQ7wYmV6t4cAX/CtOO0
JmcaueGFSzTav90ooIbGUlOv4MnRsNBBMoqGDqAlhQyQdF2I1LWoL4cjorubJpb2ohTpHkTdh+MW
yGITKo6i+/VmJSMuYaLOYs/Ak7ylMG9vuQ3QoDrGZkfUJr7kiYp+52tqZmxtSoJCCxizQpPB8TkF
Mo7obpgVg6EsTPOCCmS4lMo3+2N5Ckz2LSUOuGZTJAwIZEP0zOSQvhoJSM3tANOsnrafYIjLMgsU
KQiDS1qH5yYnanb1RD9nLRyIQAEpEiZnqlL7vkChK3ZepQqQscTylCafi+aCE5/+FBONmu8CS5bh
UZMfdK+YdfJMDGuYxvCvZP3pejjM+NahtXee739wTrFkg1gj5HOefP8LOyNvUsGKmBwEFhzkcCFZ
A5iESMBMhAA6S8oFhZQarSUSPM17nk8xD9zgdKZ4PGzOVb55zMxUE+OXgoA7kqRrEru74htNx86A
bopikA0i4urFMJ5buJv7s5f+AiJV0TdNbkhuqZU6w5E0jxxZyspqZPeIbU5S55r6sGKrFOOYUbqC
pS92QR50s8YmvZeXn9QK0mvh5gWXoLOUVkE2fo6nfFf/6W5rgradoTvfBqosCHT7nCylLSbgRXmB
38kltBU0PnskR91wc+Az4qlEDQ3EB2IcdP4tSIbHACUEmaLJ3vOT6ULRNSJ5heuZHWxV7U7Ogkqt
uYnKbOyY/LhBUnY/ZhH+fKQuiYVaKIlLONr0jy25Cf9yhdUCGhGbBZrsbM7hhsv5E6DNWk/a6Q3F
rx+NBucpG6GviPcJYPk/EVggCDq/LvF3kUma+5IFe22JwNIy6lA7BPTU2oWcbz8aV4vnCbLTcHf/
vzBmaYgtejX617Bi310ZMpWm/m2CSo0wQQsq/J8sFLlyX5TpAOpLFwGdhu/AQs3o3JwELAYW9uXr
sm/eQ2Ok5MDmUpFjtkku5Wvh5YKBRbsneAU/9/fweo/FGiJZtbEkErUbWZg5oWXw3E2rzpkM7oaV
ZgLL5Ms2YEhtFTzrJ3dyiwK7K0CX4Rly4FMt1dCfzLEDMLK8PCkAoRYocqM8DLBK9o4lKOMmtV0a
TuZL9o1ZJ1eY32JOT+EE2ykQ7G3ye+HESLIma2mtXiq8tELxH/H8KQxm4XcN1FqFFIB3q/0SBlbm
llO8eu4LiF7osh0PxgSsF/n2q2qwPYa2kIxxSVjLCjd2dM9XUO078XLadM13DQ2OiwRTQCHS1NW7
ifBwpXvVof3aU71/rYlp5gNdn8epPTtXa+i8DnnE/HfEspMWnsHhTOFog1jjyfeeNbI1EbD4pDGc
fJGzr13ARRFKG7DMp/m330rUkeq2o7vnr9GbtwEtgUctmdBMKKAkNUCzSfzHT/RtoDgWGTx1CLV9
C2nMtFDlqsgiXQ+P55O5d65xrQLk3wByM0+lTez/pXJzjT24ov8v4QKAo/x6QV5/9zbMnUIbRXzv
BPzz81ZuBFy4KrWNOLjOrUQg/x45drE9qeIZfPD5VGuO94ou/yyQlzKCQMMDYHCeU+ORWcFMVEBj
yfa4kc5oSn/wTxBSgG38a3sh0MjZhkR2t8kqcIMDDRXHG3ViPq94EIWofRANJ5R803FvMNaJuFpF
xJnpG9Ki3QfRqsMupYoWigBK1koH9mmU0bKVMm5kRxachxU1GUU4RNVznrccr/yFtGQyf6oKwe/w
/J2yzHH+3n+krShF/Em/l0567mZpqECBdXJjnq9ISeopT6CD2BuX3PLhXCnB+NQ/6M6jVEZ0ywTV
LRT9oAV98iUMQoUbPhifwGxJEpF7auVxjsQP0cdhjDDjkqH/pYEqEh0CQ2XDScC1R/xorFobeNL7
zs15Y66W2rXp+hWTi57YwK7KtWEs4fHFBGYPKtzYIEVLsyTsHzgbkUPw01eNJQrZ2JrZzuIxZfTA
tlMwT9Y4ZslaZXBFPohh5SuT5MY9jJmG+A5510uun1wukEa1wAS8u4OrTzDW/DqlmDeqbva1a0Hw
gcIik9Sjd1Rb9q2QXFh6/eYH9Rt/uOMLu8EChLVBngA/54UGA4SON1qDFeFjEInccWv3hF0vj8ly
FGwbzoO4n0a5dWjorDZqKQQVCdDIZONpFapy4GfallqAduIvOmST2slQfQSTdX7H13QQB1naFNla
0hN0R5cyoklSUNdag5wEhyK7+3ZmKr2rmd3FQMp8KZrxprL6w19t9Pu2nGsohFW6W96uNDUD1P6I
YNuCjrvWTSbvC61/jJI47pBwr9wF7ra57CCsVg7S2JA+qFV16Ci1yVY2o0MPeONyGbrCJ9GhhaiY
RYLafBvKjHe1Hviy7SU6bW1bOpBzz/SBz6fjx29NEOMIeT0oeaoHllFK+15SPGmk+tRUwL6VEPCc
7oJL1P3VTGT0AFdUDjW0TPwUVJ3mtVx9I4xwK6vdq9+obab4KoyV6rc+yAcYbvYMWzWCbzGCElxy
MPm5hN6p7XR8Di+CDRtmqMcm+7gVo65uSnPhVPaJI5lTq11s4GB+IAQpOZJMhBP+lg4ucSWdr24s
zlbiqcipX4meZMX0n6R/crnTwyFi6lxAGfuqWsL2+Yw2aNa9dq6W99/t4RwdbT2BKaNthW4hQ6DY
vWYY+mximOaFIfaCj2gOX0YFVieke9EVBehvh2zs3VVg84MP9k7A/jGM8ySr6S+xkgtasEn+j5rz
IuX/cUYsU0MIy2g7RuTp+NgbtiUOjUYejawAPCaF9s7JBBg5lYbPtzL5t5IqRwmy6iejTMkL7I0y
ILNzK4xo08xowPBfJBoWVE6eZUHyXmdcRTTSodzqPQZZOVclWkIn+Qdq7WtGv828+gM4fABoHT2y
siqQbmGFrSXyephRJ7wMrrS253rdoIr0IWeJkE/MTQSAu3Nd82tyeFZCKPhYXDOGPLtn2z1Rpejh
AdgnFbgdmc2kXiQ3HsdXXkTMygUS8+tVgM6H7o3Gomb69HKTlA3g0qANaBm/muWlWR/P/5Yt7lO1
T7fykIx9yamhtU6wjullXSzmkhAi4PT9drDbAC8rd7P/gl7eQRpaZ8urtVGqr5qhCRytzDc0wfjF
0p6gL6GJVEviJDOeSj5l4V3xlJBAeP0UeQvHOUMMOYX96/YyGMzIWftOIxvZgSWdbZZEdhOFKq5H
MNR24Xzfms6Xwp1sn3y9z0SE4fvlL87w5Uebes1vwGAzFEoe0vKnfgEPDhM5AuyLuqtWCoTeojrs
/Gmc74hjcMP1GkEq/cmPuHQ2E49Fy4+8tf5G0mooGaLf0veI30nolZUNPYeZixA7mD80o0yw6u0Q
wqn8FzxIefOfkX7KWAMObKBZTUjLr9wVPv2RAo6mKxwjJiq/8nIR+8Me3pgJ9CtlS3VtfqVgfi2P
IXKiMUmaWpD0Nuw8XVf+BKb/fLhkJytD+Q7QeOnjTOu6/SHfxPdJ78CfVda/EdoYW1RNrL0A6Awn
+pGd03YQNC5rmaHh2IjMD27k+DMMFPoxHHQSIIGO1M6dNlqyeD4LAdHxszCBO8+exLxxhbnGr59k
bTAOewqqr52En0HnbeYN8boBNVwiKPi8faLGG2HSd0/uPqKnP8EzaXWot0DuH0AOkREHD9xbvQXZ
BomDCVI4DgycbPqh+ss6xeV1kn1g4sd5rjlE8oksLwbjQ6nMY0UEVTxhjp2RzFp4RVF999TPkKwZ
UiVlXXeKt1PX91w7ZjKzFQP8kSlRaH44lNZFs9nRacXMIiB7TfnlLdOem1p3Paagd/MM0ng+HyNm
erPzKbzzbRrKY5f5gd9x0AcqyOhwKqxj9+SyiOwH/7/j/nYtxeOQqzE+r1mQpwhS6dDWzaoCQvsG
rUJoGoYt7a71mBZcjg6pc7fOzIDYKPhbU9gXSDxWVoslT0j2ZeD/ZN63AfkG3a/x9K2BcXpgybiP
pSh6zG3oxowbI/QKa+Yr0K4w4N2Td310eQOvetqWQAkaX+xQqKUG9Gp+kXpwBcWiGT5Nn1Tlr3LD
itb1wxL4Sf0qgIhMWEfg6UG7xeRW+9YSVw3uUQXgsOg5pgcXQvZkRift6QkocxnDRFtt7Xtv7Voe
a4jaFPr5Hobuvd/0CqWJklMiFvJ6JeO9Rck/OkOqc578oq8n0JAlI8MJPN6XAcfXLF8kP6E4UfmB
Og9dF6XrjOjOY3i7TKjC5Wik/nhvzvBpD4AjDUZldsvgQzRHFLXnM354Cd/YbNGFGQaeF1LppC+O
N8AJqcxb/qAGm0AZc8WRxPEcmBR0xXGbDXVWgOGEKj32j+FHs1zEeBfa2il2ETpZqefau77PZaPN
mw+VO7+ARxENYWLkq1XGYhThynL4OXRsCca3VGtZ5Gisze9AJYW8aX74idiNoDqQH6rIzo0aV4Pc
/nezzGwR2xsViC4DTTp/vtNqkE9jcMmcaZH3iafJBV+a4+ZYMf3Pkuch00F1a99JbTB5/YhYpycO
EcEV0dXFXcgwEdcBdD3moU+DMakRVpiymFNANb2B4L2HuNgGFKwrh5R9rYBUOBNJwZR3WHZwSUYF
3kv7Mc5hWCKh0YPsuDLImARJuzBGrH5S0BfGgzmSMvWmgrjBEvs9Gxt/1Q8qpbBnExlX35ZUN6Hc
IjN/3NtjhDJWvwxR719FbAMjeCRiKgek5AllwWsGiOwuKYbcNKMAAPgXEh4KH8zDY2lzBMK11loy
T4zVWYJ2wg3nidsk/m/MvcYnbYQpoI2JTbM6RH6g/TlfnWITCiwuiJZJetyxhyC19/YCucxLshA0
XcfJar3Gpnvm9NnN5EO3PLxjtdgpV5qMZ/0KHVYUjjOZhwR6Mn+URiNkdfb++jdFxNXB/rIzaNPI
s3Nf+0AQ7a86lE2zRv3M1uu/t8qyV8isoygkDt56Ka3YlA2tES//HmShmISC8vzGA1aJDl00IGvB
tejvuRh9GLukgKkb0VheqquFypXtILs662F/Ff6mx/ZlCZiZhxaEmxUbN2oVVKUGBDb1Dr1l0F9x
LFk2NnOTukhhITaByNLTq/E9W4loApHsgBblmUnxBDTSVVslY1VOhPTVExSFRFJGZuRm39cejzCg
VUCr+p4bI+smsJISt2zz5Lpi44YRPmg6R83ug6gBdGKHgOGhPQI6j5Vuz4dQXGYXhqKKgD64lCEQ
MWPxZwK7zqJ0u7DKyIMxpqoXPsa4v1g/EtSVPHGD3FR42j37WREEVmsOMpv2OshlIoGPDJAaEjY7
tCsoE30K7TN2rFFB0jj/5vH4yMX+ZMPF/durtdxWKjXSY0wfsNHK4UTUdrbWB6qKXnGNOUlDtxKP
zHlRYuk16Lo/wUikxxgQg3RNNOfKBZJD3qg3rLr7BReLX4xS+d3hGWhIhVlb1L1BKB5TfnkXTfrS
3TTG+I/oZVZGJZnf2XuIT8LR+ew8Ra3Hr/2lgpyh966hIl/c+Zynju91enluhQjiYRibf9uHE8uW
qoM2DSQSpTkc5nzKJ0Lnii1xUL2WF68K4VRJIg1KzHcZ8KLhu8mPxGSTsu1PrpTYm9jB6nMLUXBA
SDXZTFtpIUGraZ3PJm08lX/poInfoJokHEt6mvu4D1Hep2uuJEaN5SfU1Cq87znPyvP/sI4e55dv
+ZNcHA4mNDIRwXxmT+4wm+mEyl9+GUE/gzeKD1KFUP2XYYupM6ASMGf8HzqmEAY90x1rSN2LpHAN
xvOxqFSHrE0BFz/2XI12ufEE7qEsk6xxAinKGDgxF89eMGcQNWrs2xc2IYlUn6lS9wRzMEqmOPdc
aTSFlZVPyEjpmCgDT06Fpcp4lKzdkE49pQhTtANyUk5+2+VOskh+vjVUgygO6uVrF3H0T0Fdg2f5
ANcBGchg4zBTl14vzUJAZLLVpjWLvTtcs18a615HqlJSRAGgp3MDJbvWhSSfxj1+EMJPop2IntiX
ktxeeaDBzS1j7Ev7yigDwdoJYOlMG3+8V6QTueCbJTd/d/KouhuPeKUb+z0U3N3ltHWiWbklXJgV
A56Oq4q38gwkHz5uYuFSWvwfP7HRuo+rPSFOoi91MD5LKqP30++3+xPnfLEh5Wl6wy06LnQ6NTRO
7a5KRlrc+tkiybei5GFATQawX6p4FWu990lkhjfoX9MVS1BdGa1qIDHSTiqsCcPBhcdeNbE7bxsC
Nuj1axq2+Rh0zSRGtlsxpXK72TRAhBeFsXLUoJw3/yWaEYGrtdxqYTDbGFZ8hV8F84L33EXcmuMt
9D/xJO1TOX3D3+wzxAWiEh2EWnGuEm6Tn2r3T3+gEwdyvTp9Sv0w4MtGqe7L5FY/goFU1DqjsDsj
OWxguEWyedwh/mUxn5GeUM48SRI6uR3v4GbnwNzu+Qka3jUHBgjMETzvFz0xJuxHpGpCGM9bfecb
GxaQ4EJrSyDdb6UIX9xhMVPEJCmUbNcFpobSYgVHEbs/ey1aiI8HN1G+7z3dG6W8ZwNxd2DRO8z9
B0nI8yExH4Tb9lxDq1QVPTr6h/dHa49/EsNBBXJn35n886v1qHjc966Z1a73yeA1AbCQS7AoTSnK
OFJkmd6KH9G8Pc82vPqI/Dz2gq92spZloB/CGVRRwm/u2P8+ssRNWK+IBC6QIKu9tS4Y8sKWmmny
hO7thCoVzO0rdkXsnXfTdXMJcViRlxdX3lmjuaPNAQpDNNl0A2jiloEDy3gLOmD0Bm5hQ8+3hZ/E
Zvi2psZB7rQitMtYhn8371+pvHoC0OcoNc4diLA1VxzfsZ7x3GUWzd9PeTIYnH1kslDKYg0vXNxD
lQ6uxIPBGH+r9EUX7W9P+is48iDdd5NAqEkzEzik5h2TGjAExIs/K5n7H/Dv/51f0RVD6Uw/7l6y
xYuICnt8aa7C28SVCylhhzIQkUjauuI3EJN/ZWMXRZ+GW/S6Ho+JupcULNLP+zFpFkwONPFCKGAA
D7e5Q9VcsAwi+NIL0RvtUsOx7nzIz3M5Arzj0Jj+6w23lvzHPi/YIPmaoSXk3JmTDFnAi2Mmrq4s
l8JwzvTZdmqcwOk7HYanmlBt6DsbL7l0rZsUIY8MZ0YPqePb24LlUOYUS95YhjzLdbeW8pc+Ep3b
8sL3mPHPgZdxpIdAHb1d6QdITNX8ENuk++HpA2p4M1c9HXGcpIUUaaM/fMjjq6/ofHu10UOJFavx
g1BshU8kp9jsGBy0dCDdwov+DiV2lhG52/XGbFYqxGMV8jiiUN40Xrv6Mu/103/Cqprwpjo2B6W/
3o9bLeDYqX9nQ01VlWZAj+jU+8sDWKyjuPhyRK84fdyaIMURVE5kuj1ttWmFROwqBVAYYfx1K+VS
Q6V6EK3vZ+VoqYBijNAzJYclnv3ctPIVUv+8Clb1mq1qqyE56x67a5XdcBsZikbYE+CkYFUprmXR
ar+ooEu7WyUq6eERpIr7hXrlBJKMcFFGQPgvCo9yv3ZgNhTe47umyrwQLoyNcGSolU+j7FmuYmFx
H0FoEFOt9IbAKaLJxGiKRfHO66JiHrN3kKMpBHnoZAaaN8xsu21rx3Soj4HsN0oAnmk0uD1lBXpJ
fvG38hxiiCh/Cdb56EeKACmfvCqVsk9qbe6wIiZYZA5SMabwdyW7gpFrvZJ+RZ8z4I421gZf6DS3
JMJ4rJIaSVlnfGBqncsiGg7v/ysijI9PGTXBBvAV+iP3PHkoyj9lBJlJrxAfHD/WCH83OMnmuoJ4
0iCKRJt80LkVz3IC8biIyzhT7eVUINRQIp6WRe6Gt3ViO3VHv/u+/76cryZUNSG3SkAfOtZhKHrC
vKhbckHK2+CZOjc3XLrKYD3mMoIgPsZdMOmY5HbZ2+SynBh8xXhDhqmzCiErzpWZX8MZaIDxJYmE
vLMuAzOmfBLV+qyfgdF2A7q/NBGS/fC7wCz4hl3XgBvBbFyaPdRyILkyoEnURP117AELywFxOzOM
WWBFIDw/MXkTd6e6u+rnmiYhV8XimVpOPHAbmXy5OercTVy4Rp1AFaqGZa55WzQf7w6e7XJKPeOt
/unXjrFh6I0J3p5GE1xH0HicXExrpBC150TTlp4ll4QeOwkZWD/25SkJhkKkSrxkYZ5QSk2NQuE6
UewHYNh7pa3uB7bhQoEXf8mTh4CfP6A8zTcEj6J/A6cSQJcELkar0zydjtCDX4YMOd3ZeHKvl5q8
EY1xROLLqvGCSO9k2Iq3waHjZhAXiBdLxLnsaVYryE3kzmvLjNQ0if8mxTdLUVHbh3poOgBhscha
3z5wDTekMiFOct3jmiV87hgpkTLlXw/XgL5NEWTKFskL3K1bbwmHOP8ovCd9ocDTHfI1TKGtHM98
+nkekNGpO2JzdEgNSbe9yjrZpXLOP/64hjUpLGhdcEpYKhDMzuIZ2EqFkeWGpnhYA3Jq4ySwjvan
z9xZQZKvLbtRQN2JLHherGTpqypbvLyLt+QvAODjC/HOaWcnd9W48iSNXyP8ZKKYARNPGJ66Yp75
V9d3cc3wtKJ01pzx+HnFO4GMBOQ/I5E5EcwZg1v7U//xu+BjGL3bxZiVpZJWM/wd+AIbc4wEbMEw
jH3jgXdxQNJ1CIy3LyJjWzaoX3c/7P0jFOGyWpMvaYqV/zO7RphnODBh/YHg2NA2UljZFTLGZimB
wWFORIri+iTGHOjlk0Rw6yzM/A8PouRohWsqUiT9L2T74fNRzCmqTqYRzxXCTnunxyjRImZjINoP
PgpT6pr8B3hFyu1RQp2HAO6vpYWJRczM68+lZPFMjMTQ/bDH2IdbKCIomkktqvevXhARmvnz5FuI
pwslIaxA0UGWsLIRZoN+AUd3BAkCmJTiq1XYAWBSAzyKHPNVRrxN+zPAO4hPgABNntxM83yKWllR
lMdm/BejzswvJjmbBnfdbaDGVoJVmG0jVHtQx7oTii5GJfpHlz+z3bPMEeZ/kyKgBZAkCIKRAR2B
K9tAMCGLgyjFQT6Fo9IYfl1J/TTFo556me4w8rm4trnuBTpcPvHB35dAvVhOj0kKkdNIYO/aeirK
git2N5fqMSScCMcPRXXuHKnrrW/saXVzdQTgaNdOxW4CJUIdCZKwuvNm/84/qWGJ2v6Udx7zv/LG
8i7HINVFF7VuqDwuUlCkpGrNu0ehjVOC0YWJMWc9m3sOi7r7qF4N5iHrqxqDBnanGEi3Lpm/dtdM
bcOtSCIVgCHOjHZwUWBGLdOHtr0RAmoP9yK2YbpPRfwTOpUdOPutTPD9DAozHPUeG/EoQmee9AOu
xg0uF/Y/ygodd4Ts2V3ap9+cOB/VTueCphUwPi2XCTG6kPT9ZJhtW+2uXuXXKybJBxyjN0uDLSu5
VAm4Ucg+zGKFSNmiZeEJkzr64G4ENNTgToLOeK6V+oyR7so4oHRE7XM0iaMHFT9Kjz01FOLnpMY9
UdMtJU4e027WsNtiVVUsXC4enAftsGGFQjLrVMX7KPQY9OmHyAJp0Dyyw7OxTUbBrr3juw1euReC
1NJqzDdFU1N2Bes0n3MoAbGnioI0a2WtaP8Ps1aHCIeacWH2aJNnIUJbcJtHK05wxvjy2zDoXruX
/oE8PBAmkr1UHXAF0tlZ5QSbdAKVMCl5H2PYU1l3u7EXD9U3sCbuHyFnVuQlc7xfeZUXf6J0vmpm
Tk1a7fw6u+wHnGa9Fdvv0sTHrUaudEXZ7oGCegzkbIiSBGtFqYpLTY1+rD8X1a/GoGvRzA/7vxHn
WcAbXSVg9Q9wt09UMDMPm/tBytxqoiYRz60Wp9L/qkahzW8ZfZuQmQFotJh5tlzxOv0gMBjVOLVC
5J89lK8Hfh60y4coQLP0ZaDq94KCZj6UelhWW80ygUJ74tAulENt9NWdMMzFcBKFsX/MqnKqc+Ty
pbKNH9dsm4bRjGsbGjsfkJZOPeKeX/GlOGWg5HroA5mbG9r/LHASPPxFZdqwM4IpsbgU0rQ62qh2
hmn7879Ws0rHznaZ6jKRMKUy+gXqVEHBfDbmZOkmEpzdWvW6rMXbTd9YKGicLggKft+eLIw2QlwB
ngKj1Gd+M5fL8RbSaslvwjrOjKyc+Bdkq0zwik2Qrfw0xCyeZVuqFIZdwcz8fWxy1E1MDMOyVVX0
YS9CapzqHbL9UZFlVDNNZCLbaAxjkkX9F/DoMK5TZXpXn70J04cMYxL4513HakdhgvIrvHRU1ist
1HKtmC4I8d4PY97fkGII7oPOGXeFLQPN+5qe95FtF94FbE9pWsQeoD+8cOUR85QK2i6kqLlFI9lK
wyrK9EV+neMgz7uab7mzV3tSLoK3ppFKiZpZh8iOOxbQWuaogJRx3WnlrqAFerjYw99xsQE1iGtj
0oo9VGYNgc+ay6sTM4L+BBREOG8JxGHvZKt36ws2bCqb4I0F/nXdzB1UYod0O7+PSYYAJHnvjk0y
TB2KEIMKLz/bG8JcOAKaKBNTYJW2OGQGYm6cgEEaWKWGQ1hpt/4X9oTgYAY+stxw+CySuy4MdK2t
FwL3+kn9iA6kEwjbCxkwNoVIbEQbL17s+0maUKBLjm2ClMjt7F8qfuaAOGDOJ3kRVZFAP+nTXG8Y
iFk/V8fauc07U9E+a/9o4DT8N4V6QJJx4lReA9TDvW4NzwVAFAxziUQTNo2H009Z/sLEyO/mPqf0
wFDtAgcjCxdi2qlPeV41kfPZn5Ka/Zy8jKIUZVE6gdifjN7rTdhBZ/VXIOhYHKIluUqr72acP19v
JvyfjDTV2UJ5Fg5008rorMY6DTX4+VxbBshpq8aFAi+uhPVMGOjDy/1eBXsxPGC8LpMH3Ju7+Zbu
wCpBWOAFg09ill6zpwK7uYSoCTxLDyb09MJa79B4gHexZfbLTPqtiQzCmCL7nVKps/5zkz89Qstk
viWoFD9K/d47388OW2Yf8qazTIoI1//lsTcIlZr5R4wKqQM8NhrXrPqd0AaNt4seu5qURw0LNsvw
RJXimPEAFrN2iZXJLDNcFT+4sudLISnObhUdDR2WSg8VgPm+IbboIKyvKn7KaQo52X8q+haUdcy5
UE06TQIbseJ5NNaK2HFPFKaOO8s3bUK4obt8k544LLir02S53ctDO8xkot+uF+FWPMYNiiJ2HY8z
ccG6Uk4JXQXJev12XeIJhqPHyQ/Oh3Tnb8+3F+QLSQ+DPphjBA5jbYVIziTQsiG1J6AdWKbC2rgJ
qrPbU7OVK4SMdrvPjFoJ9ZZT1H5dnHd8AV3Ahfmt8SPcPiA2uGYB0qg8VsEg4P/Q/hQSTN9Au185
qyWixGipxPXhArU10C4pwgrGdOeaXotKKjF/lWhqZWUcWw9U3hUvuwPwQGmLA57i30xcA50ib4+V
XEtPG+VezUCctirCXHeuPlGQh948iUrT92JDyouqnzVS7JZQdZg8PazXsBJ0XEODM8vqOXrwuP+n
uGrcca2lQxVqaY4dQnhppKTdndG/ta0W3Qp32EAWs35+VtPErPsXGdswE3GSMeU0Ao/ySzrdOral
U2AL6XMJcJGKv8FqezfWjS8nXIvygbKVqFixaQS6Wr1X1hzdpOa6fRN5TAP/apG6ztY0iGAZb1r0
Dj6KwgG3J85icSmYd2AJbnD0GFgX/eRolK2irgG5JlV1F8KkD8aRFqPGLQJUJxqkjzFOX4irAUeM
FNR6eZTiJIObO5Sho1+sWvFEYq8Ou5BmSAWQKo0l+Oq2V9BKnklrdco3JSrzNv2McGybKGfReOEu
IzsYH5eHqGsgXyMl/XQ8RCgkmp4p/woCmESaUX+Ji6sez8ym9ZMBGv6g2NMiHUs4Lx+6tDQfykRV
ZYCEE8Tl0XyCCaYvdp6yKklmEjABLxpZv7cm6e9Rq9/t4IQCR9Y1APueoLgKe+5UUnmS5+12FMss
AiHFU2r3cR+e2f+5r/2bcSwd+HWXajTiouyEict7qOG1y7QWffh2CwxN+YtlzLtkAfxw2wlh4edB
WCsl6NzIJ5m2WnYr990xJJpA8ixT/030UPQDZOp7AuRuGgWb5vZF9nn475gS3Sj9O0CykielJlTe
M169qAI4DdeHYdvMl9kkPZte5lWm77EnoAe7/iM0mZ5OQejIqvfd677C+JMMP9+YvUI6XGUKhDj8
Xmb0S9jk+DsLJJE5qPjg18nO27ucbASpfeTK07S4y11yyf1Op+sBR1tx3dlKNTZYSOZf45ZN8ver
PLoY2sjbVQnBhmKQjN+R1gUIj8W9o+2l3CLjoSM9fCGqhI/123BG4uGsP8GJkygO3TZ4Uu3see/b
aiH1EPYIQyfVFymn662edxh0Rd8XOFyDZw2ndNt7WEXt2rXSXIcNz63GtI0eK17kEwQeM64+el/r
BjiydonVZbZ/pdLrkosqXznsB85ApbcpaeiGxQApxa6H0SVHInBRGKDugqkV6zOuSF+YK9ZSIYCC
yzXb3IlUSoVD8mWY0qDzLOo22X/eS3/Fh7XeOoukY6p1ZoENXq6EzPY/ez2Zr5/vBuefB5LSdA+V
bYzMklQ8MJykEJ5l1BzJjl1IuBdLRcLTxI1UWI46NmKSe83H/DWEPUraXQx07jqH0jiZuhrjv6e/
iAPJcW+LJe2ObZSaceTeN4DXBR8vTyXVPFQ3ZkuPm8JIhhuxY8iTCVDZxDNjowb1dpIzwb3FgQUj
s1WZiMNhMwltNo83nCe46RR8lEI7m4FjPZc8hY+oO0pYQrH66qBYFnO3nxPlE1Pvh7ZUKAE/V+NP
N63xcfhXxatnyrTxBkbbavSCcsMoj0oXbkq8Bllz9xAG6NKzNVRP28v7jiyWW1skrWAGdh8oo5Ya
ILOjCaMk0TzM44tp3jDywWcrBCj5qut4KIq2F5zaShJyp1PA0VMYl3wQwJUD20HFOX32Hi9a64Q5
Ojr4sATECn9Byv51JpM4S2tOSkKn+VoTn1b+Omw1kstUGwQaBSWuoyCRd+75u7Bu4aU4+Ts/5L7/
IXIou3QUnv14KoZ3/bKApK/0sgveE7Z89rk2+M3qUNWfqj+Bof9tQ+qqiD2Zk+CjEOiczK9b50ov
igDqtC0lzUJMM41epQ2t/wZk89COO8yfKyeQLHdE+CQGz3kIxrtaAxCirFI88EkM/d1CU3lqWMWU
NbpQNcRTekVIvRymXn0TV2DQejyq41/PKWm2a+WKbaE9ZrS3BS+aDp4PJvBf4BMbLfkYvBUkfF1O
V5vNi7Q7uVLeY8MPo253TE+0tvLgDvh6UJlkN65/FyeZUsr87Px9Bi4vxx3vssxmp73jBoM9wGtd
AMGmX1JKq26ArW71ThE5O2YxltG7DyqcJG0OyDOFXOm4Dy2aM7Q36kYoqWfknxXzsbji5+0ckqZp
Qc6Ika6L5z7nI8WF9w3Z8VFL02ih38MA4RCl0QXwZcZgpxouSeA97MOGU2JCUtR93qYmsReja13P
jyw7SxmgGRVzxHy+qkf8VYdFOzprYm7g5lcB9JdOPYPFQmpRtK2zoSggrfnOrIvLhm6BWG9YXIvH
svztDZjmxaC7EMCbv8qMhDMYz2lBfU9dnz17WsdB7yUJ53CC7AuyfPDEikIY9iGwAuZgGhBymcDM
nrmCMVS5N/htU55ByKORBCrUqCAQCVWPrLlgIIEsRz433rGrPnH2jcwMhqFIvtfpT/Gux9cZJDIV
DW5gGOgK3NqfiybtwuKVP2r8XNA1rL/Apr4Vl6zubVbyW0E9KM0exSOzk640xE9V09UKwgm+zzUG
hTKxO7fqmQilS24DiEu9K0Wnvb5eogJq683EtnlhOkvLZI7y6rVhmmkzSZCDGR7MR7RtFpk/ezF9
EL2j4YJUltJCKFToC3tFyJLncR0PmCPeKpG3TZJs840gk/xVRXCuSdDL8Skgb+jvoRNigrkPN8q1
QURUj16zq90QnqwmtPa9iF+e5rdil6Evhn3Z3x70Z/pgXcJz5Vxf39qb4DuUEizFfxoMNOcMKeEF
6PJD0SrywKhgpo0u1vEdKnaoHWjUgtHXzW+TvVSpI/HjVszKFcJC5CQjucaBsWOIi73oF57daCOV
z/cq3BFPxBtTOSyz5CgPr55BlFhXBtrEapm236YEgeqkXxhK0terM59klYXD+CSsJZtidjZfidBq
2u823VcJdO4M5OFlVdPQUJXiThQGK15RJiAUBQMBbZmIfH+xxONzuO4YOnB/T5J/y7bkHFX7cY7z
N3pgGIxK7Fn41aa/LFypfepglxbdAU0SwmPFlsU8m4uQ/i2OaLDye2U2Bp/kTF/51WU5Zh5NENZK
TIhjUYoIPCndbqjzHRGugCtvBKVSlgk5JvIkOdg3Pf7i2CsLLY7vKhylJg+9TbHqCsJWauEuAkul
ju4foRsUdCmHVR0oLj8WpkQIAG1QLRQTCYo0sTFwnygYuxs5g+uRdSuAZ/lyx9wfXnIN8M1keI2u
ZVagK4v8bxboJTrZuppZm+0TRZmxcHiZUxz8fzZ90XV0acpTy/nFBGkOOxGBGVNz5oZv2mxXeCGF
Rh6l/+mvEt76WdqMFcRcvnR/DWwF37hvNI6Is3tDROzWjqtab96OvI1RDtsJNXYcQJ2gjqUrn4TC
CLwhLXIX0X1ynCko5ZGVVjFUIX5grsx5eBNLGr3zlG9n7hqu+lO5kDCJzuqqB+/DdmjfD6Ilsbfe
VDfhHrVr37BDN5+B6WpqVzT/PAu4ymAPzDohbEsB3rbqSw8i5ThgwEi6iYMoZYQueIZHJqwyA4Qt
AFEdo052OauwA2OQJKLrB1U5xvOqsM+4i+AjSFMznJYuPgluo40eUIic55lyqADSI7UJSUNLQj0F
ivfqYfjK9Ne1iEa4y63OuM+ZLVxKOnb8/SxIgLF5hOvINUuKAQ+qBR/b2QGLCGki+pthcvrGZLvn
728l0HU2PVTSJN9h9RZX6itOotghIVWEVCkbfqaBLHyc63Slf40gadO/OXMRVcvzLIvkKUL2+GnN
J0A1dCTGhLgaV2ceq0nFOH3hwafo6h7Y4v695/rD10cqega1UZFXsLd+UvP7W3ZR3hqdclTlEkYI
+QgdLvLmeDfPrHmaP1BhwXcKqkObafH6J29Dd5khDW2FYDmpKOtGUn6ojX6PQs/g/Rpz+7mA0pzI
7TrEc7MGdX1sMMlmG2BU0Tm95agA5S8OvPka0e9F+Xsc7snEaOkWnVP0ipIzc9HIQi16IkcoxJbG
fxXcg/Y8daPeW3k5SOed1qdVRzauJCMXGMzf/8jd4ax+1DEDwX9Mso87+sXsemUUtLdj6OIp21/F
ANNE8Tkd/kr+mjQSPr664HYBiWx2N42VrTSIzpJo4tI3fQz+2etK4D0wKkC1+mcgsjSr8AJhfKka
Y2tTFvqUpk1aMk8AzZPruhUBPSjcr82mEZ4RQImGpGwRcIOeHfDPlCrEVIfGH5PcV5u9o1cvH8gK
JP8g4k195XbOBKlO0BW/F2wNKEzmkEkiLzicw2a3U5aJzSy7srKh1b1UavLtc5oq2hW4dTaruV2p
eZz/ege6DQqXomPHzYrqGewXri6UcGjLs0Aa/Su7V3D/3ctilJ0sgxqIGnsItRD+HzT+9ogELbK7
D/toORARKpJc0A+St//6+p3rEwiW7K7f9Hb2SH3uu7BoR4vdw2/FZV9AsfpsliPY2U3r2Vt69tdn
M0fzYvtvyQdNnpkKogv7D3r1+bgZKvFWQ4FiQqv/u+l7uDxuutQBwCHjO/diLCbUwNEuUBbBWoIO
XzIrs/P+CODD+ECWC0uEbcdwBrQOrZAu1+QRoLZDJom9+3mVVKuZOTub7MPGUPBgFa9MhLv93LoH
VdjRG15bckCPlNYh1OBkUveHQC0bTqdui0/zz1xOtx1WFkDlbv7PG261cisOifXPJzWpVKOH0qYq
WyyK+plpoId+KnSRM0wGNsMZ5vvXFjkuPTJB7vdgqI6g++9iuYLCe+e0lQUi/zecy6OvISq5Jfnb
BICQi4L+3OJ1Ju7aZ7BFT9LfKCUFo/t4lMwkjbxDGdoBT5tmynVjkzHILl6aOxFbrItsOM6sY8oP
xO5jDyA2lowu8STx0kCNv1lHdrNg70J6ZjulDhKq4FOYJElvageKxw22S2GzExM3e48Dnqybgw3i
p7XZd35DZ8utv6peQNfmiGOxjkHKGXwkDgSzVOXTFoyUN8WxNP1MaCeFqfPNIz5P9hjFU2EQn+2X
gHpZ0raiEEkxxv8c3kqT/cGyhhv8kEj2GmnCSFIEk5bk577YzipgY18CCnr1ODMmoTLX022Ir78x
M7Q3Vrk1SQSNeSt5G1KQJKs0zxva04Tv7yIMEXYkvACvgHZlvNV68JZh0RN46cJGO9G8fqlkcnhe
SnGBaCBZ7pDoCPBHKN6B/ymCM7n6W78WAlOvDn7uzPGOf5i1bNc2cB58comppO3yY0VKrmR8CnDN
CCyrUbE9mDP4rgGWPUkMqBFOgTocDjF7utGiW2KUB2PqdoXXeDroEZuJhUj2An//yNLIBDTPbRH0
F6ZzOitGD0tyOo9PGE8w7/svnwQWyyv4LNmM2kEWV7gtlOEU6rOs9dKLod5pkmiF+Sq55JeJv7Tn
KQAN2xUsq9d5eusw7GUbJcZwjQFsZHo2SKZePvT7B+jcYgEsmi3XXUovahJffyn550/2c9OJtGAA
p7eNNPRrcO9lauleuJwT2XunsGYTpzst0/ROLGqfi7GM7U/DqKxAwX1XY35Bl1L7SgYPL5dvw8zA
kqGaAm0YXHkptPON//BwB4oZzdv4MM979kJ74qt9Dz+UmWQEtVoAQxw56duNNZo9lfmgOWirfWSg
75Us74aciBSq+hUi+kmUMtCs2kIY4JcF9Ev49la/BfMGJY9ESvDsKhr4eycjzd3kuc2rfZ90XFFS
YkLAdFtl9qoGvBa0lPxR0p8GCrkoS6r3WjPNRXsCLs7CyXSv5plyj9nyuArHTtf8r2/YAhglmYdz
A5hpOPW1lev1de79Ad2kAK9V3+FUti13DOEWrfBkZQXZ0TPWOd2bJKXIsd8/fqg2p86mmcy2/701
C7daxfaUJlwytHakfvx4KfBuAcxv9lPBP87aXne2hgJGV2jy69I1y7ZE+Ztx4k+NSk4tCV42YXmx
5WudHcr+jBfOCGAMjL2x6LAezGrCW6hRF/w30NxqwqMqIBR1X6U8H/ADoU3fCQdgjbVuZQx9fzpF
aprUY4EcsBBEHqPW5QD+9BDhVz3pnnPIN4GXy0GdD+L0Z9DoEm3lflLo82gF10sLmNOjaGUU7GiL
OgO+cvtWoqdPzCqWsKpCSdeQEF/CJ4+6q6tEQQuOlXN9hLwTltF7T5AP0CK6ExVwhuwFbAlJaRth
RuijC/7VlYitgKuwXgs1kU+PA4Lzmje1pxb1XHdmX7EUTlSpjvDzr8d3JEdkSvuJm1bzu9wEi8Br
KUSZQc8WnS7b8jEu7h3VlAJdtXl+Z8rGVe4d+SMU0pAwA57H5jeiEJFVZc5E0tU7HoLkY/UyqGEs
J40sZpEx5wIKxxwRN3MZub59JfA5fQ5U9+TxL+cDBaozProm4hTRclj1KNrUCWhAM6+5upjq+JJj
9gSxa0t9tBv1U8bPCX+GIyz9PiakNKu7u38CE3MB7I0Z8XxHjzJu02sVY0EAqtR9gmHP33wBWQ01
us4okKQJ0rLV80EUvb5OLQyxUVI7spdfpKa8MFCXRByIlbGP2dpP4eElLzAOFTu+WrihElw/Rtk+
+PE3utjwSTzNL2cUKq/qw3StOY9MmxX+P904azddiIjPXplvKlM9mbuu1VdnkEw2v5y2kD4g1DIW
LmK2LsJ3CyPIccOwF0p+Od9NyxKRMrOEoSqX0kFGOu54Pgr0lahmKku3rg5smXv1x3I6htkgf2p5
J/6HBNg5rIPUGnzBr2oYuAjaoePIdKGw7XXUKycj8cavysTLbwseIbn9W434fA6HcbIlvRZHFFJP
W+dzX//T/qYtF+1sxwuk6MXs8gV2/rhqFA3Wcrs5mT/vGCvyx1jVCySgY8abFkf5+ooF74nCyx5o
w0TrVy2XmLRXI+b4dfpofjjY8o3h6o7ZKt+AtNLcbp/x5Si7+bv0uW5cNuQUlfCpVAhxDE6SNKEm
lkAxSFKLIHUsFwM5Zrt6SLZKpvers9H8BRAnVznCeDYCcuDSsX3q94FlrCvrvtfA3OM7P2BQVnrf
Hrb4muy3tTy3oWows25p+9IcIJheIFyfhmGHpJgt6CS96CZDgM8jgJcZvK4AxGxp8nj7sj8LAY7F
wVnBCKzh+OIVaRsjA45d7MltEIhYInOsCpihIiL0RKfeuY1VcCYqUz6soOVMkrmj3Bvg/jdLCVVa
pUlmILf4Yl44dUIRJjHNmq2sPJTP3Elw7xhPiy44A/kzMM6JuoIP3n++NsFmbQt+8tiPN2JEv+/E
i4u3T9HWJ3NIPuep0qV+MMLVeZslvRs2LZUWOu6PpsgSqO3J2ENA+5WCKDJNtvvM3YD1ay5ViYJp
BqOIvwBNEMjusL1plk+XYT/gqm0Ehf8/eh7Byo62GyAg5XLaa7mXNMOOTMFsgX79ukq4iLpi5QJS
/QqbEfdSH3Ao4/Uvml/Wsk44FVWyLOfB/lEq7YoZ8vm5bty0fh2wmUOlVqlX1mc7MRuYygw5RC7q
IQpXRyKa412M2IfsMsJm1poLRCKQJDbZB5ILh71ScpExivTexf33dcUMQC2REkA/uC2naaxmFujt
jOyeOFt8i/60muCX34Bpr9YdsY2aIR5QgaM9bFlDpkCqMBk1qnxwuXIr62pORL10kNqOeEflCpzC
PkD0vcX8hHvm4l0RZrIM4+QisecwQHNw8U45S+z41SOt0+k2ceKjA48XU2V4XNsEvyyfdwAe+HTl
KXXnBxRFUSIWiX+8ty52l98m7OyRQygEpeUNQPJCw8aV0bWmHqdT72Zb+8QlEAiYKOLpHcqR/DYM
QGrCIRkTerwWtgNKemHlnxNgNzuO4Fmm3cNUoLSrYYPncrYdseeluy3uTLIdvGLcUHfC6ZCaGGlA
P50/RH3YV1YncaVVOJTIlza/O2/bgFtcusiatf+pEDOQa9NDk2nvNCDGH2uBlrwO4oGnn00OE89t
H4jmDPXrILy/zx1CRis6BukEMf1lDjd6jVpD0TkZaVrEpM/HiE3JIoiT4OYjdPwNEpwM3SBfksGa
QprG/YORrNCOacArLs117G+v9GSlXAGzO9Z9dZxQ1vQ+FKkaC431Bl55GqLTFpXsIrRIf0K0hlR1
plBYK7hjQAVa5CVa/74l0fGB6yQk1/YWGYv77iNaklFA9l+TuslT2c6A7cZQedfKXitgm/4Nkyuo
jcrPY0zx+nY4fWIhElboagSQoy2uXOjcH2XG7KD1PE+GRHnIMi5X7M4rgBamzfr4WabLdC8tIqKR
3TATdRE51ZbY87ZIEx1YRqFcjctV4mc/dQuudyPB9NDB2j+mtk19YXwZaZM0H8/p6rwuCoNTG7dn
1kwSC7BAWwt2W5NT5n6G8uk5sYEwAQ9pI1zCxD0CQdhxFqZsx+asK5CHEYhlqJte3uFJ1IZElTlx
Fu9jK73fYxf3rcR9mJxOWakMq0m9H+mAyjKKvevO8sxVAaLDhm8dHpYy/KTDsSHKZITSuixI1v/I
/+NZwPPSb5lQOIvXNxmYLRpfpUQdaIlyhVWaSReoVbR2tz0OBwCrm6snraOFv1r37MzI5TmuroHm
9ft5hYU8KWzeW2Lsk6p+Apb/vkcK5YlM0l6b/twK0cO724+aejVxDaxsLgCAPkeX69W8BdU/oTH6
oC6hlcFwDe1rHVNqlva4MJcKo7i0YZ575DcaGfDPo5q78NFpoLj0WP2z/8gbNWa+4V26pvo8c3ix
O4X3g1CI3/Sw38oW15zTjPqVA7SuzZOZKwDuuSAHB5qBUbxHU2espWTQp5otax6LXCoywrHgafbT
bwA8ZSXtVYgrwtOrroSWIRgoXlmYaVuQcvtq1agdU/968IWZq4Plhk/tSkvSYExBc+gL/pcDG7FF
5jahEIkERI6HVo3urO+aCsblyyGy29puqrS5MyRXnQ4nLFuUvbJ2qF5TZhWkpsalHdmiBpybrN6K
WZkqH7MSvoawtp7NtObrcfypdfxhkp4v4B2IYL8ABRYfMiCJmKJmbDbvVqPvuBE5rLmoojgR7UZq
DH4ixYIgmZlQnQuDhF/tUZyEDy6yEohOfIgAXeKnIbFBgLl+Iua2Nh++Uq8S0gRd6qO9tLYwhmSa
w4C6G/NZhqPmhIGP3gij/LZKf1353so57nq3szNPm3KDzm0/oJgDGdyXHV9RzyOyyt7j3zzFXuFN
77q5pujORWgikncw2kDADCzDNuFzMgmiJY/O/HN7hwh3qsjqX+zQGU42aD7PzmzmCORTDezAg4zZ
q0Kk7NP6I+tqtOTCG2BFNGarXG5W1joXLdfAUL/rud8eh2P/J8AnTZc7pCvYgIrYMqpP1H9E8cP/
lLqcEvuYjYL8PMcvDr+roavKt3zL7TXhg9f9m4Di4PcNGBHxJbRHgcXyZC6OlZeQB+dPHFvmR8qi
dsA0sr6nvdBxJk5s/GumiyRMmoATYbZwgQHL6ok2Xy+YG6P7YKhvMRC+gCyE7SjcpXR03b0Ujujz
R1SLsdzy73pL1v2e76WY8JTgeLJUw2xMorq+HuGe3LH0hZtVVy8TWf5D1S0XtGcDMDCh9zTU+i0E
iO9qNGzFA3RYae5avZm/RplUN6YrysTl3TdKenuQEr3Xk344vvkc45e9Mou7jViOwhgZJt4/AFjW
r4G9Fu9W4ddWVWlCW2o+sYjPWZ6lgr5eMFWPGEMjqxzUsUhHO6W4tSBx13ZB4xHqV6A35NLEzmk4
4QjttIH8/7of9jKgMi8zJGXP4vwaR1DF5dewodHPk+oqJy02B1HWYukJn3G8SqbJ3ZPdZQYYP/Cw
XlqkNsTBFxcwCvrpaE/e104DaSkaalyTon3/Nx+IgYcOsFCJU6H+fQO+qywrkbPhRKYzT/4=
`protect end_protected
