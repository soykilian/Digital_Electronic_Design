`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BzuWO1rJgaA0PGodEZCyhHs4oFdRklp3Tn0lwa19mhVB5ODlIC4JEi9GLqZ+EMA440stL1QxXAwR
phcbxabC0w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a+x6i6LfQdTq6YEsKd/J7ZCNpm8z+SLyk42JFplkMCCqfOIizSj7bdU+FsZRXn/iIAt519f168Zy
sCfZLq0o9O8YSNtfIZjCYYLMRR+N2r3wQUTorzdf2/NZdVjY5UBMtpsSAlhqlq/kai1RH0/Z5Wts
yRK9RefQH3rIE+6PncQ=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ex4YSsJ0FXhvUfhveSyt+dWXJuKU63a5ugYfjLe116Zc+McbHrbgWTat0Grt9eDVmRVxImMKucbd
z10CElrDq0A6EA+HfDoSekW8Bi+2UwvVfBqjKGBWlCRC4NXak8RcIwTs67M1ZdZWQRpl3yja0phc
pEdMRXCNG+2nhGcwnBk=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pwPdjPXC8aJytre8XZN2fK+Sc7UwXBKYK3xU09qGyohDNc4r9MBfLHcBEriH36fL61VXydQnDRgw
z55n+IfgHTePwdZC/wCFQfNEBJ9nNbj5xfJ8kz9oHnS0DwSALXVOFonc512YUpl2uOupJ6FPED5V
DKmDNxWGhuF1hMnw3zNrKYX6ouqA5K0UxD+leGpbHD8Yt2yO4cvRff0/u+PxA1CeJDDwhgmsxS3V
xbCL4paRo5smveLwGDKGxyfCrUlIE2hssVXFu49KgGWEJqMEh/ZeSjiF/4pMUeamWfXrMFE5b0lS
42CPUwoVV31ktb9HeJKDSvBdG8a21Z+VWhd74Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HklfsDWvQXqz7VjMwDP54j0MK/CyXnBIHjFSVzYwt5RmcFxEbVx1CKjEf8Vn0MJk+ogX7q/bVBut
iHRBFggKO+h8p0k2+hClN+VOv3f6fjVlSs4lBSqokAapvNsrkpGB9h/HdY4kBLNpZS2uPiw4z6yj
SXq//+UU4gZBUxADQNtCb+azWQHNnruF+ff9cQ5j/ZDcfqPOmjiMz7aMuSWvv2fBEmJj+PnnSjNK
bpNhtVSHqARpOwTXE+EFvO1+mTCJ37+dBX6FVgG8JPYUTjXkQcpKjmf+cnGXkC3sSf9KmLlRu3K9
sCRoQKUF3ooA08pdnFcB10MtZgg6t2N14E/9bw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IRi2KjPb1F9FLQe8XAg112d7VZnWdwpc1p4VMKUXFC+O6s8GyJ4xzET+82u7fXwQ9KiRT/C2ohU0
IKzZFJ/VgCo/VKel9v8rgYEbHpZ1N2HI+yNDuC/Gpxn4Ny8PAFR1sCqvmcXmM4YkvOpEPjTGlNbQ
OfzkR+0WfGpd1WXacmtny0PQPE3VYprBWh/NwUDWS954TEh542CGmGePsCyWIJhdw3k+8LBj3a9B
QIbM0vS8KOMlyvY02+daccN13z3hMnqrssyC3bW4D/4FAhr6FvnQOhr9unzZCBcVwLcDENauA8jQ
AOJCtvAutMkASfyeY0w5o5g0ddktSDrqnAl+cA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 121856)
`protect data_block
LqYTBrc4Xt8HNs56IUnEzx2BhxefZNspqxHxvJ+zrwZ4SdVB5gHxltCXlNizfMbpPW9+Yn68RrfN
U/5I4+byKB6cIz8WKWufG5UaX6M0ij52Am+TRaGR9eqmRGPbNIfqkCFXm2LnWJlaCyxa9R88vWcx
cPvb/hWGrNNeYS86OGwu4u3vpN806ICNFgkSFlXXv2+i6nClP+e4DBQxOy1iyyrji2NZybXi3TZH
Q3dveIKP4kwZA4i+mUhBlXKTVvu97R3AUX7csNofVmalFQ5j4WRSNjHGolbZoY0uGgREMT99EH2s
lr9+ySoOPCwaf6R5WQ3hsRgYaim027xgILk7rP8u+qUs1U4Nqd2tH7ZJy25pzDcr3gSOS+zTdMi+
TBcIKGlwT7AC2kY9oUdMGrZwfbIuBZfK9/EHjibGAuRjui/7ZHEzoK3ESSgbUbQWHpCoJi8J/ygy
MrazPPo4Hw+eG+ZcivQORMS0phqwOaU53GUlDcoyc0rW6h3PE4kjkpTbGMUjzFCejKNoA/onrgB1
ZPr3PiCVScPecotU0hVfaLc99fGZjJsKIKcf5szNzUgJ/FFx2KKYJN4n7CVe24ZC/OtYWZjhNCQa
aTcExHgaiQMuuT6ZThHgIGp/H9T+yopcc/ou7AWnVZyFj2mpwajiYf3DEpRVMUYiVm2udF+XECFD
ACimkRydV8fZK7xH7+CX5GZMMCZSVVtPrFAiFQwZiYdkH1SnW5RaZ5qeHMLbCVA4OR8kdb38b7Fh
zxfsi/Co3CLn06BaOy/ckUzzeO2Bi0EBXFVELATpy/DaPcjvMOM19iNzwJc3Zle/vvNQfqcUg2Zy
+hlYJLq+6xTbCaq8RpDr5GV4THrLIVU0FMq8RgYMBOqROT2DuhG4KPx5JAGCiBRgG8yzygqbkcWq
Cn5Ub4cNGA+buzdMfcglIsuHi3g0dluPUmhVuUNQyN60wNY1riPFtZmBW0mrFfUgxS5RKRhsJ9ai
25MjyxYFvPsHAql1xFZHcR5Gh1/1IuXPKXPn92HA6zChVgkSrK+EB459tOC8iihyS8OjSs+IcEbw
5/fXxAi6Xl5ERV0nN7zaUzO/5Kwl+Svu7+flcaA9JxZXI9VMwNMjkqLc4UxB0VVdp/YgtJ+Eeyyq
tK1ZkVC7JH7Fcxw0SO2XWtZzipn7bTol51MgRVbx988recBHCaLbhoCSHDYwD3SdtdgrkRm6ottq
eN39vStw/unUw3orexcUowT/LxtBD8QuFHWqQz7IoUfSH9u6WVsw6KPVHo/Pj+m/r+qiyKv6rNKI
URRFUzX24vqrTVW0jQxgGVkdY3WptXQA18+uqiZtayy2gpfOYYvKP67NJZGtH4wpkxwXNhKvy2j6
7wBDr3e35WT7tQnYR871cih8Y4cZF0mBY79oiPN87irT7CnxpzAKdB7VEuH8k4lt56jhZ7F6mDlv
cvB92OLWO8dW4DS18pDbkabPs2R5faMk1/5L4yaklKyo0r5hCdIXxSYoVGehaa0QdAT4Vb1znWrP
dhOzEsFzUUwjl0yvGJruZugO+gCUjyB/kb9Me4dFh2qWugYiNCPW495ukA5UUxM0qXSaSJSfOwd+
bjHRET0KwRIdATncqf2AKv/xmyQW4mDqp971wH5C5PhNqv0ZGNn19n0TAYSCcgWRBR07heZsODJq
Py1kO88wAnUthHgncIrfOfjSda+Ata1X7lgQ39etmr+ksbcBpt6jRf/beHQIbw6w8LfUy1u16uYx
H7vGY/a3dNIOY7QwJhKFomL8seDqjCn75GOO7QYjd23oVVSFgEtfH8DjCkUCK42hn6QmNIw2QYTp
3rdBxczBVlffY6kFZZdbgYrZk4SbqdvNa1CPiCrJx6PyV39qu3z1PuSpFLzUEwKqA8B5i1xd5TVr
9/Yo57bc10tuG3tEUeraT1GFbROlWH47x4g9mp8BvccLKwfH0VR2E7MTkd0T8fQsDx+rlYQZ7NFs
5q5PML5Q5pAummNzaWjnI8d7qse1gvIrxrRF9W2boU4dsKqc8nlNyXA9SSsvE0u+OQFrICRpiWPc
d39qHdxMQw7J6D+PY0PNiTAWfVAAxgA6QaWoOGP7W+Xxb6CqR/sSFEhO6LCmpGWhK3+TneS8Dj20
X+y+c3tP7co4nccLgU5waDktUT0IcSsdmNQmNEew8LI9ZnQcP3IFGys6819B9GPq4Jayzwo+IEg4
c8LlBRPFNZVQjlMoSGv8uTzNryuu1VUzJHycG+8SGNwxF3BkZEr1+jBZqC77T7dr2PXa+jt6Ty0F
TCuQ+HxAI0KqWFJe46/aZF5LskKl6EbgI887iOcJQcuVm1GbjLHMUsmfOLQZCy3ZnYBu8Bl9VZEJ
7ry1Q7lzsBTpK/ZywxED9pDME5M/dhQOMUC3LPGesS/9qZ4xJMBvV6z6O6V2B9kMtVcBXBJNYgzP
oVgYsmMmlH9aN9PD2CNwXOxsdrqrFQvG7kpKaz4dESKkUxiz/wG7w4CKmWR9jy0XYr/1qUq48GzX
K+zNSSRKE7SvpKvYchd0F/E6mLd5+1bRJe6EHCJVDNhQF6fiaTD25wLCG0xSjrCyZuNCQ2mATkcU
MgYW3IbIVeXp9A/A9+rnRICsd9fXnBJG2E/KfaA8QB2tWw1S6bz2YmXTznOJFfolVkVP4Exn5rQY
TIlZxSegcVLsA2Pm5WS9M3zdarw+fQamikIvB/rNjEUtJUSF5zKbNrPxWUKfj3On82mK9Id51t9G
TrvBxIXAPLTVQaP3sOxIo6FC9QQPcItaDOkJa2bW+kXAtmQPaPcDqQdeMCw/ORtHvBlPElzStqnb
xZTmHp7dVUziu7DOyzIVla/52ldjQC0UVzBnaoIJzdi7ch+gn32pDShcMQM5FGaxzBQQRYLT+9n/
T+sgSq+Wb2zsfCpJPOzEZtIB+5bF6EwFEJYiGgiarJTlBokzEa5Zoqms6hsIPqRmdvGDzUbe0ioK
abQG5Ay7BSy5loG7xKnrgmMKEP2H4be+CI9jczKTLbukWoVyXmQnp7hsyoM1vBF/whjHdAlBAMBK
9hmVOGrpoqsC9hEjRY4S+CWCcXmB3mwXsTSvTIOSgDKDc04Q3B4RcF+XkkjC4i90b11laNiEHhUg
QxHmAOD3F9nIU0WS6MO8XAd6LJxv1vBhTf7UHAAqdXRtkvp7Y/+fJNWxe2/F7aEWg8G4qyu4+1rh
SB+m+ByDsCmAG8EBpJvK/go/Ae9H7LS509JAaINB4s49ZHk1ohDI5cnz39qcMs0tTmFvsD0GgpC6
d1bfkb6aGcngUsxCo9JvGSzYG8rvYLm7r5us6BzgAQJvuZmMU3D4zbmT5vm3gYhv242fAV9/5kcU
HnMWgPRCSqu8QiOwtCGi1qW9dowd+4Iy4XBQ0FEk22InE/O8yi5CEjUvXni+AFsaBFtMVqI+XRni
cRlj3QvgkWrmRkRdVczodZnSKEgC27olvgHAuUHw/EwrqBN9CZIik54LINZcaovGy033rryNP4w6
uctXjRJAaEneO6YJurnVYPraC2JgUB/NLGOs013c4L+5FaUVVvb4pKNtc03GuNTrtm5s8XNhHU9d
W2pkF5iICk1oGecDRWN2f1H4esCIQE3ba2q3aBXUeEZd56FtSA3bGaBX0uB+5fh5LY8sghYnAoiO
sX4Y3/JXOCluKEQuwaK/xRwE8uhLAEc1f1E32JxH7XkpzgSdQarTkYiOcekae9kGnz5Epp9MkwKI
kBsA3MxYyJwBY6YT2VmPcBM6f1QfcQUd8WdQea0R8dojXx4Gzqyn6ukyTLzETX4nA5nrbKkDFTRA
EUbqOAHRj5RljeKMGiRXfxu4+zd1U5iwvKFTAVLHd5KyO4ocKLC6s4ys1QGbO/Qac3PlY0AXIqo9
lu/i6ySZeqDlmo5tfvmMNkdT8WhXkKyddgtkkXjCBlDL06kDi+z7RGZQWXZoCUTln7baJau3xX18
oSF4lqyx+gN3jtZEmeRjMEOEgGRz/VwqfymwBTAEvLw9Vv8AAvZgzOpYIivvIgQlMFYg6wtQ09It
RkvPPvRW5hPzPw/fWwrRAk+t5orFnGpz8YQNzc7XFml0xqju5hw3e9lKo2XK2h167BlXrdlBQW0g
YZdPg6sZ/GGCM+F8LGvX0cn6XUFnfa/CC+rWSwuosf0X8l38keiZyXnQHWaFeajJ1rO8unFdnKnt
NHxhQ3uNGJMbf+oI5IcunS/EhWgBkIBF1VL8B+X6bN0NKaBHk72cyy5ptm/LjA3B4X3bFCQk2ouV
HYUxkpZxCzyhqunhzCs7fafrXDC41WOdnBebhCS9Z6DZ/TdXJN+ubchUoDpNT9LhvlwLLQA1aVhJ
WbkMok7curlIcSshqNaMkFvYc5LhLdFqtydvVBBfgXcJMd4hD3dUmniGc87wjEivvuEL2Adxo7yF
a6wVhq908lxNDjzwSTjKHW+it9Ts7zR6b+0tTN2bUZSX9CDgBNIvxZ+nbW7w2X+yPgRAjH1QZcbp
eGPQF1FlXBSruQXpS0JcftZUcGqAgO274Ja6CkRtBOFRL0pxJCxdIQzNA6d+73b1hnpKBWFPdctn
dA4pOjbKy5Oc58OcSeRJ62dBeROWkwwJh2NoEFeNjAMFQYdXrl8qiKWCT1rQdp5lqhmizUwMRPBW
1C7EjYJHgynn2Va1YduQFSS0bZRwuYphnzKU/mo1z/Xb3yJYNucr9k6JOdAiwjZ9q6jbmwBwMLqn
p9iwWKy6kphIZ2xAsnItP1vAFFAEHPMZ1CtW/JFVXwSCkiWGE8R8b7k372x1IzGNODpRRxFxPMMC
OS9haiohPoKw6eentuG/FrAYtosbaSrISimtV4rKJfMP2vFO3+knVpHfIl1RwASrq0KATIbKOJtr
jFkmvJErNaFEh2thy6hni8bfLIipxcz1P+HZyyxCLasfpfd3MZrdIEpMB9SyiuafbvVjxwwagKrc
Js4SFWG/1fL1TAc+jyffuPwrko2FXoWOyshpyIH5sj4qh78YRa8q5ssz8HjLU4sCoZj4a7En1Tqs
deCoE61Re4CXmOsyBNsDnXVFBMR0JEyiycg410oi+sk3SdOCOh81PiPOp/1LPbeSwBiZpZcdxoNd
5ff72YpRO7uUSxRAYovUD0pzdYBfC9CUiVeo+J+OrePRFJGuTyDGpiVqzVDDiJyiD02zPOmA2ZaW
fNUcHd85isPEXJ6ObJpDOAL4/DzwYBfMwS4dnVnjyQApSypUsWPHQ9xv9wcftCkHpbzayL3LbCTF
wMQNKtXm5BHr9+3gTapkZCOBcQVrY+rdfeR5F7t3TVJXhsnU1VaT3q2Fnbb5tgUfJTSRzoqsqkoj
LH8bf7m7o5ljXPO6RA7pgWb8OPJIIo/AlBDQzefD6kzXXjV54JpXEZMoUMh8DMEOUP/B2aUh+KqJ
pzD3x7iYJuGzIquOLKeMovqrq4YKUc3X8w9lAEz5GLCtH8U3LRxlRMlolFaioXIkBwpWJXg+731r
d4xmWglK6093CHlD0OpyZuRT8JOnZc37iZIl7vPSUOWNe+whcWrr61cTFu2iPSma30JnZGWbTgUU
QEClFu8HB1Qy1ImAEd7m5O2ceJRdZLggCxesiu6crPzhYs8wnynyslzUav+KuuMVgiXA34ffDvxq
zNkQ3mAu+hqESAMh+70nXqwdEe+q1lA06iyLS8IcJfEmK55CwNxsPIG6jFPQK4BZsjF9PIXi4Ned
1KppEFBRZ5k3dKUet+k3rMyEut5OPsROKokxKPKx9VNIfYx20y0NCXdTKe2oPfUlqkBlR4po12ZK
yK9UlT5rvcF2zFMHimFFzia91A8B99NX/32yZc/+wKKZn02A3TXSqExrHTgbXX8P3oumrwP3F+ga
scq1y96szjPEHbBgtY7DGrfcpeDpE0d88HdXziM73oBaILC4yADdttTV4qPFHcPL5juhsanw877p
sXLH+HmM7WfYrkDyGNwsHesbYgi+YQ29RzSHXBYmdREc710bEIi88AGzUSgE03/vjRBL7EYfK7Y4
QrrKNqmnXdCG3VzspAyPgVTmJn7WrrdZFfwZXsa4dHE+jm8obGAKU1eztg4SaocHeXggLZmn0aO/
SWjr5+SLTqxWSeyBm6wLS+HwgYC18orZ5j6cB24Brjs0WBoKB09p8gJR9rhnzkiAo/kjxS7GUUt/
YuXfgHwCDgMCXRPlYy+JMHhrnA6fqihWQtJdpqiVKyfOK1zu0juwKLB+ZYhKKIPQSqRTJmur8wqE
po7bbcGt1s3EGhYSIYmMOyS/7XhdmsGZPqSTQf3u93gBYUnjpU5FlACbfoiOON16yXJN1SL5tI/o
2WerhHFbBSR5VJgL1sQoHBJDn5mRfBQv8ZBcppddEVwS9gwZqGZ23Csa2vTm+eYn+t00ZNXM76af
OJ14A7Xm5TlH5+ZGZagZu/dqAtXzr8LhvjgKkZ3RxE6m5OqdIbqvPimlZrP2ylBPMJg3bW+XRp1A
dkQ9tNEgb9mKLfk/B7B64g3cocJ2N5w+vqSIZfXUvriVKsjCvCc0KKI7RbNXITzCKjwkDYoeUvzT
IjWfy+tW3/cLXUIOmTR28hBVquZmPqb1jut4EqeeULkgOFhGndqmS6B0qcWJ+EOe1baJb2FvkDCc
TuweRnjdvz88ay87MvJhCXpQHVzioWMHZfWMXSF5Qu6LIgECcYcGvvPgP5cIeez06JFHQXyFVU7r
fdlP/LD//AWZjjp95TETerHOLBd4HhadzRl1fPvtU25zcNEw1lkrbx2dQ1+N76KqypT6jS0sMxAe
z3y/iQen0kmi5Pw2r5MGEaxoggezIepnlSq5syIlboKzUrSHhm4u3UWeOhEkq/wa6Iyd5yXsrHao
35Z0QkHO0H73NG88MqWmE/EslW4nxvSkhbV271heey5k8w2U8NN3wYFo/pDu/3LU0D/AI8DMcOlG
hLbEENVJMoBMWwXK7DgvnJUFr9NhmmuHgJkMBIT4vRO/Yu8ZijUIcLtT3r5DWVP5+g2koGMcrSLh
lgXX3j4yC1XeLs2iv14BipwSvfL9RCOJD5p/EoTVWKKUoz/hvimO7z0ydifTmrq9wMeoq3cV9XMx
xlPcKySb8ZFzIzyNt7ls984jx1r68drn8BRxgCPXHaJdKb6pBMbacDtH3Xr0ViAHXCoypaHy0yGb
ycYvJfVIysykvphdvKyQbJXVd6J8yVoNrxr45GIra37B19qL2sDx5K4hZBJh6wxsk/tmraXUYPB+
79vmNQ24bH3RoiOOnfNaDIcAOQDZ/PzLP6EGK+ABMNgiI7w1egd/tJO2+tLmuuRJBMrOQhsIaAxc
so57Ist+X4vULhjaf+schnZQ9aFFLBRouXvNreEQ2V2EQb0QAjPiHm6fSrc5cZHUdG1y4H3Cs3kP
g1SnV2JIS6PEFrEOBl8aeZ6SyLnro4PgDkmCEfIGsVynBBkJwfn0a740e9VuK80Z+6SJrWkxcGaV
iXI4C0hxwBmqfc9wr3MsBv5bElINNAvZGwtandCaLMGDh8TuiW0VrFajrtuOYPrn2Y/9Z85FEuRw
XW7PGCEOv300yjTUECHinmtbPC7fg9KzBerr/tPEWEeiAxQtUbbGcSoRRsOFHZEkXPlBh5nH67VU
Iu/l/GgTGzyl1sNfxRfvkf3oiQUL0QJykext+pg6S1Xi9YL7C7Gnq4nsaAC4YJxo8WSowPPWQqOS
127+YSeq8Mta+G9szbsWCXTQc7MK0QISiFf8gu24eV6G3asrU8v6p5RASA7zodiCwHHGYrJ/RlgH
nOhrPw8YAn5nVPfY6BiA0kym+zc5TGQ2NITmANILI+RZ0ZTe8SkPpc1J7UeFwcyH6iM34c3OwtRA
qLFIJGoOyvnzJbrgRpkj4poEwoSjqQQDFA7qzG/D2K3JFQoV0ghjtstQaIN6b5gj3Zjg18XnkMuv
7dr5clFUXDObHHNZPY05mkbTCtRy2C0EE9aeqIkUL3sOD4/kpWzhDexx88CYoENQ8xLbJP3RIArv
aOdjcJZMUodgr2ZI2dJ0MwNaWJe3r77AqOLsaTF1M7piUM/PeYjExSgAmW518aC3IMRKFFy+1OEV
dHtqEhsw/ibfizM1OaBFx63M4EoAt10/cRLy6fGqTJIwr6WM0rHFdPIAJwFa8d185P0K0aDzLJND
/+hsnitYM6yZBxOMs6WRM0MjLnPkxLRakPdz1N9ypMSs4mTXwLLHt1qiBGkP+KZag0NjPn89occR
Mmu30xI9J7ZVrVQn+H83yKbaRzOcuVFOdYbhNamKIEsP0ff/BF6qTCal/sUbfAAou8ikFL+QzLNi
GCuf587bfmyrRk/CnICuOqvwYh00tg1YjmQCFiW7iopqEfdBnDaiRc1pbpX56yOfgNEb4xGqzKr1
Df1QF0oausLA7E5d6S+quw8INuYByQry1qQcZTYAsMSN2/Gyn1k3OGu/stQTp6EEthikLPnOoeb5
USYZBfPpSGA9IWts7S/PK1zB9hGzTznhFVGjsDsxTXoemNpFZnhIEwdfywlCZp0WRvSQfdqFsj5K
HWUXszgeSCT+pztobaJfbNM37NMJfh85rDAEVKT8pmYYAYcQcJFzJ4dDT85bqURdjZtFfXWpjQ/p
kAel1Rzw9LKfJW+wGBAQh6k8X3qf/so8/NhIBMqdJ8ZmcWGyTMEnzV7tqpt+wbTOnnW+dbu8MzsU
hApzrq5d68MUC9RwHhZscd4jhJ/I/KkXP19eXwIBXBDIs0UNmBrVxqADDx9OcSmlpaT4iIjaYXLP
+KOgoGpEqSOTdnCXAtwmCJovpedDi/5ZFx2ptfshsYi7/ZiXPT3l2aGIRhCSWq3rOanG3u4RFaIP
pGKjiNTmT+TkJzLCZsshlIes42LuUgnVv9REiTnGhD7y3vawW0QRothIcqpKBTyN4HnW9vHVb4ea
t+wqtDfAof1YHa61wms2XEpW7S8iI1ayqTK5wNC5WT+2HdBoz21rfPpNfPLKI3vwAfoUN+jeUiaQ
ElkzuU5O6795jkzT03GXg2usL/LTG5r+6/0/CjsTzDXnWsv21qhjMJeJebZZcyshsiP4IKHa/q8L
3aFJ06zsliXDZUpdlHgplBwP2DsMf+2cijuMcgjNFqqhn0Dc1RoGvAjPdTRu3mrEA6Y2rtS3v2cH
89EXzmEnoCRLAtQoqBwMu296RYrCD0i+5rzyKDwJYI5TpRYWDJCKkTYnJXomI1Mtqnfm9H2lO/oY
aiF4Vo/DSOO+PuxbboLg8aVd4Nx6DecxbhqUpJIMFKNPkRDb9LbMCRhHINed5UmuE6L0P1YjjNai
oXGof1UgyyNd/a8Os/X6SM74SGBVDRFKm5Qxiv2KwNkmUlDaHYwe/f/Tt3Nrmyf7tfhMO17QLfQe
iOrnKiNqqzePPyLZwR+NopCDQbktdwH1zuRLwjQX1O9oTKrSwPB0zCDBWsGnKlvQ1snoNGEwdCxW
KSOCFn7tCmXgRNtpKHXvB/YHWwVLFX/FjxpxkkC79tAOAFE7up6lHPFS01QRm5N4Qa0nFJ4lBSaO
Fn3JUZTaVKvRgFbmkdz132AqaVYsI3z8cX2S5haNCjATHjRSu4W350Jdc5jQcEA+PtXI8iqADSyb
lK57NyfPdV5dFedUwMoZawXUZ5t9RscpNpk6LDklhgXz1uZsSfydozhU0rBDtP8I63ghZ51HhwrQ
AUuqXq4h9J0qKtfAz2qIRZXF44X36f9VMcbkdqlZ4Jvrc0e0920XSexYDi7mISroP6MN7Jn5EEaM
KQ+IIkn/Xz3LYMZf+dO6ubSw/5ruajw/WyFtDbyBfVl7CBeB6+1dfA7puhtT22OECDMdBntRCpvN
B0ueG83c49eqB/Ei2uDFsZJ3xQEgIRwteX9+x4IVEzoLcy/IfL9ZBbrfSV5YzZleWTMU8D3SCavE
ZaZ1yLrgt9029DpOQC6L//3Xqk2bE3tlYl1SatjJKCyRRmFSUykhOu7GfxWanKI0x0V4elfQiPfg
H/QXl9N+8QYr7z1gqdTGQ9jPSJH/Pw1JEY8H7CZa8wryCdG6IsXxODYMxxE+xfEFkPrbccrHrjYP
zFFLMcB/2AwGCtab/qS++26ZWHBUAix00UTtDTP5KS6luipBpsdEtuCxaCq90cA282dK+bxz6H+9
m6BRUbGCdVxOPJVYu+F7yW/W3MoNTvxbDeUTaCauYmGhP626N8q5QrixfyqjsxVMW9d+LlTzDzC4
HgCJxAKLXy/W1XAi5E4nU+SfPZEAFUJ+dYChuz/bdPdpys4sQZQKVqLe/mcBke4/Pyq2/DTGF07D
q9PVxoPrBPWomWCAzs32prSzbITIRAJvvi4S5Eny7cInjKqA/M7Ws6AFlfUcf2EWeE3uRh5s7rB+
xuiiLrIBd2tiJyjTBLpBUSlfMRi33ckibf/7jD7naf5OycgESd/i8d9E8Sx3/GqEauFwq5Lv8fF+
fGpwqMATT0Z5fwXa+zuEsRyJiLSSc6dk3xp8bONA4xiYCxOJS1PeH56Uv9AqzaYdOte6WGhl/R5d
geGeiCyJ0RB/TdWsEEnqhTkAQ/v5Y8wMcPkFuqtrvZBLrBwEmG7vOc864FgUJnzTRAPXBu6Uni5B
4m3B5vip2O9k8FPNQ0jFqmauHThKfOBZPhH2i62C0ZMFZbzwnNRL2EteQhCyaxveq7mGzLVg9XO9
sRtVgvIRN0em2A5e8UYYqFDqP4MZ5SiA0CdFunnyerNNERA/ktjKTSfruL+dAS9sSVWwIjdA87pc
mDq4e50qR+tMxFD7DcMKZ+AUVNcUklEwTZWncwY2oOLUMqJvZqF+N5C9ulzGfn1Vsi4s6w1k/PFO
5n9Z6mE2dLWxdUlRIadhVTVfTdGrsHUo+ncZR7a6yj45Uku80KlZaR1U4mXZMCuP47CMIM5fhBlb
EPh4crACiu4cMl48i8ZQQzdnle7ifswX5z+39Tbu3CF8VK8OFITVtqBkyd2r3MshsuJhluTlzf4Y
EM4Qm6+7Q6jseU90pWjQmUS7HRCEBFqDh5lSU2yHgUp+haFqq5M9t8WsD0sZixDUDTBEQmyIcDJG
nOSTha2zAApCQKuyU/KfRad0+L/JXFbuNMPACXZJDKYrui7kuxU2N0H9sGRg3dzrhExRhRnqQKOz
wJOl5AHAnM2sXSVQWy0Q4IvpaSJlORgKf1PasWed4xS+EKhQUbj0QSPmOW7EkLd9ULBYc0mttl8k
NTM+0BSH27LitbfOC+3DsSvMq8U+/KmijJ7L/sNchvUHCOuylUcoYjMuZFJmDcjBpMzmvbmiBRX+
oDx8CBYC+uFOqwu4bsEhBg99kbQmprznv/pPFGhkbyB370FpY5/Gk8TmMcXlTNOQUH4ZWnxsiuIQ
2PYJaMFYy4tTTe8Va+6wrHOOGAL8YIi5tat36I4f240qfk2DFEkS5m0+Ny6EpBdBMvuPthDN01Y2
enYhf2pPi0rdEo5tfdrURLlMjoCdr6FAoqemYWev/4TYxukwMbR28t4iFO1QPJ5skhguc/HorOPE
BIGKQ/lV8WgMmnOdqMH1cHss4yWQRNSySXrW44OvNESojrxn4rBQ26oULAntAmienUcgVcY+cuhO
jD/4vDMQcyHRZ//q7obawY+psBeSxTX0EMxzi1zseofJll2oBBwp0nO9mrtNwapaMHaot1NKMnA/
4EgCy89nqEUjO5MQHW89cfgsYafmWsruswbDwISzW08LciDCJDiCPSzg2TY2eU+j4umvJwTb6ikJ
Rpe8ccRJM5RzzHGj0FRClwVl9LbojvxyR0hRy7kqX9FJWMTmGodGwYfYX94V8JidMN+k/gBBWPUb
xMS3Hy2A8lPGSB4nvhgyckcMDKqxLBJLhA7OASMtWFq1hIztxFLD/zQfMCpHjeqiqraEyzOhr3gZ
XggvAMGbbWYMopC8MpdYza9E1Jh78Jag8uoyy6lTLLWNJd/9gYmknXF9j6eb4FE10SfCSdsmEoGd
3uHdk70DMUTbLZjHjfW2BLdn2p+ZY1IiYGcL+FmaIkVI+7p8bFN3ozJu+OV4NGdr/+ajffTYt/Ow
zj79fKXxQbK5NPfpTcFJhfSpKNG6tYCI3O/nSbuFPpJzncUjhTetFaV+Iwn3XJlXJfWG7Sw++MAX
zk0NaU3z16Z+Hii6emPB/ilkHJSzyl6gDuPAkaqYdIdXkunLdZAahqjC/9n/OSiVlUnl9lUW4IrZ
Vd2vujimaJUSA11VpaA0ubyrSeG4L5YtjkCXwy3vFz9s4ablR9sEzPOJztX53NZnpZnyzO1lC+bv
iGC5olFoi6dG2sapcg0k4aKF/OfSGW6iNECHWy4BQ5jcQXM5cvmr/kP39MHdErnOpb/yiMod1EoS
9flHA7HCCYp/GO+WsosU+DYs+jxfpGk+wMfNhqenULiYt/r4HDU4WqvFKTW8KBldaimf0EgYz023
QAC4ZRiTyYxfwRXZiaaEjjHSnPqBGu+Sl68AZ4R6JAiQW9j/riibLRKsPPoPhWtP/9sderKJWnxX
kJfBgxg2VeugIKwcKeUFwoxZGaDp5uJNWsAdecE76AQiuKBxwmAc5r6JAGgxwJGmyv5pjZMcivPQ
O3NSSQ2+XLv19xE71c5JXvJZTS2gljeDxyZ5lsO/nx1iafWg2OHDZl+MZ5umW0iDH7sE9Uvqmw9X
U+rR8G62zfaTpt882yTZJB4xKuqtQ22LOIs7XWpgVGioXDP3gBmm5N0UeHjPkR7mSJCVmg2MkYZ8
zponiC5z58fOgWpiHih71FC1xN0py+YPFvrakTy5OKVeEqDifSHtb/R8IGOTEGmm0yrd113AkMzP
3JEC5dA0dKGh2a69BaGPvHMdTTy6atTizII7vgzR2lhiBTgb5E5lKP6W2ON7tOmq1Nhn/DlFt9ce
2orUDPHlokD2l0o2Mn89SfBweOUrBiu/7FyuUf+Chj9clvHJ+gjT8RuixX5Q4cjYi8bpYAt4qaNO
xUmojGpNfeAhotdRLVhxjMQDnz6Q7x3vTj1vk1JEIYKD2Qe7/NdwMcaBkdtHoyV7cfJdeQGJm3W9
Oot+o2ds0XCN8XMKQeT5dIDmr9gW25yQ6MhaAz5zUMKBbtnWXJnaap2Bff7c83280+h9dvvUmAgp
YQGWxlbMyHs+1/zRff/YD9aZH9pjQB+EXvuhUZuHBtrSaYsxCsW6pr20BQjxLCm7Am73reK8VRMm
GWuaPrs0U4ImxkMEKxs6NAveKHvk9SP2Lok6yCyBGlX0xBHpeoq7W+jDWr37Te+mQj3uqvr7zXhM
DCta64JQ0gB5yucA90aKM495Ab+UfMKwn3WcgQDnvJ+VN1DvD57AkQdCwUEUw1nH83IzbIBpSepo
4XYjawxaLqWmJD53pb34Q7mU1XyfVapOI7dOBkS52qfCsQtvCoVMy5lpEqyzzJoZ0pBdXAG4DQn5
MMZJOPs0cfNsAuY9t8sD1IljrQn/dnvYPHycBrlIvh5rAJS7o4MnFupDl93w1h9xatilZORUY6Ef
+6m7nMlDUoe+ARurz1Yw1uS0NTE6jVw6rrqVca2kN58qY/wKgI+4jfQKf2BAADbXu7j8LsciVJRN
7Q8BUocDO8RbfpfeKFR2MVnQHCBG/b2yBZPci6rV2aqC9cL0TkPaG4WxJQf8T3iyWUZ4QmwFsm91
j0D3cyLrRo0YIzyPjg4XpKlXY5S8d3ZQ5qkBDmftHAkU4tvHugTLdCVvRa+LBJiX+UceXv6l5g8o
K+FcXJbvJVFpXXV7rVsdGd4J3wS/BdBgUcFz5iCwDZejwP6QOIL3IFAYbw+IakEEYKHSmU8+pUGH
lGjf+2xDdpU+J5McELOsKPHwHQF3ENSMGdjRJwwcSYL5biQqjmVR9QJivNoyt4kMR80KAa0yNhvf
87AjCRL3ukajftFPVQWQkZgQyhjMpMaFqW6hQiV9niWqpbeQxo8A8FVXxoQqYpd1DFdeRNyqFvEX
isexKKaOmLcdRDhptG9l64/9SbeOwMHazkLyCZN1Q00g3JRfcqV8vO+rf8ueQbyLVusfPF1+nCt1
KR3AUYa7/ACSZmVtN/ej0QdCNvsrm0ncDc6lRctge+WjjDE3gjbE6gDSDl5+ek5eD+V6rwDCePTS
wzDIqz6bilIzZEsjNmTpZFaGL4HfsFIvnJImL+y3IfwN4SEnAUfJpYHPyfZX4v+5pJPj9XZWL7Ls
nE+/MvzpAl1yFT89DhmVwMUKXNKlLjDew9BOEr5WrlM9HQsO1IPcJFd+f58Ujpmp2IDVlSK4nMJt
9p3wJsySOBpZng63pS1xF+2/UAktQlT8EIGsgJV9LwYdYXF/otHoUQK9x5QbDByyIDSqO1u+hQ6d
j242NneyDEtAtok1nWwv5osuVGhGHh+lBlSo4oQ+/IoXAZnzx/K7GRk3zxW9JDyBuCg/o/qEAKVz
beBBsnDBtkG+pRk8VRLgmsvwEVHODcud65ETvHIRQ0rGUBa2F44E/k2SCkkBb9xsqWmmIBOteVyY
6Var+rCA4H+bBvSSSOimituF5ZML1yC4Lw6i3eFkt+zGCJ90xIy+aKOkEU7xjjli2rjC0z2/yevk
ZBs7pztYPIs9XKQB4LSJBaWZb3Y5EibU/SqkhkOp511jXLGCd26wk5LAAbpa8dU5WGxqA4poHNs1
O2bdxErRqjmaTs9KL5WPxebfqEgOi9Ly53IyYO93vSEDG7+SBl1WeoBDoEncB2hV0YlnQIce18nN
Ewlu1QAsShSJh71R2xXkMMO/vMZ+kiJpaLZ6l7F7AFyskBHSObaWO5qwnPeTT6Y/INUn6BTAhjUn
SQ59jo4WwduwVXWPatY9jYMPwzyxlM6vr+ws2MlpxRVn+CkpehrXMWDpIG8NnV/8J2L+j50gnRNp
n6K7m8YIKrjbEeoyEg2azdCqi9yUv3mUyULap+rq3RjOjZgR7CS1rx61E7zxxvlb7wNveiPASohv
/RP1FzxUR9cceBw6jrqHG2ADQataoRQ2F9ZcfJ1V4qMTvJ4tZMiTKspXE8oypjHQiri/DuaT5l+F
rxh8OZByDTBDUagFy1QuMyJq/azQFwVNxm4pxy0PFR1/zAp7RB2hOhBPEn1ptJRI0JuJ04zFETCv
6twr+O4A4vCmFN/OtujtyhULr0CZ7M2bff4bkhD06tBPmfFMWBNpugFN/Qmpk0GKud4JAQJe5Fdr
wemP2wyCEC2KLvujvOxhSKB/8rMhwDgXOdH0zw+JeIp77Wj4jcMCY0RsbjOe/SqsFXg/IU8TRt+q
oJdOCicBaFoHB9Ta3bHBbsZqr6nHb6GWgXXqKbywoY5zhGNy3C5WN2IdUVoJnGTY4QNjr3I+zfL5
lJ457vIqbkBBDb++BJmFVpPXa1pfc19YjFfMGeswNo9RysJEjJMwwe0w1A9yxFAANijY1F27AMMe
YFXQvAS1ZKUmWroom3xKMrhEOotLgAB+vg1Ov2p0QyhFO+cG3Zid8iow7UgSu/GUPU74kt4Ms+AZ
AoXjT1RDat2ZlQjzbQeQlhj7IYI5mZ0/2Ty0GmAELzj7SMWWEEk5fpYdmP1hygAl8wMKvO/CVT/T
Pxf6NJTvfCopRKqqV2/6uWXBUL+pyEYoxtSCwmVw2iTd8QwqZUpxk4lsGgJ4uhob1rKIuAEgz0Ca
ltSlYD3xmZFMykMZqCl0FC1xKYz/9R2G4h1zZ6GDF0voZYOkBqfA7m58eIrAu+M+wP4STiVKqcSh
iKa2hU81oFuyIh1HEVcYMxXT5BCISSOqwE+O78WlzaYR19XMlj2HtLYf3WTjcX/9uwDnGf5JJknk
ijA+rjDD2cvMwGy34uH7/IQ54LW46pBax9/kE8aHRHmNprs6uOQ8SYFLSopEyFDGcuTSFszws68v
GYnSdOYLyFJYNLjrjzYTH8VtQYj/Sq4eui74n5WIvwchywj3zAwuCWqSblZlzNATH2MSrpT6bX9q
jSs1Suy3ccFw8hsFoJ4VTTdh2aiKzkf8vSKPvMOcofQ63r+zUaQZ01M0skePwvfn6+xdc95Iaf5Z
OJtva6wVLTICkz6X6lI1NsWjciOu6Tc3CrFZvvtfgoj8kHUpRyjLnO9yQ71r2iwl2gUQt3uWJeLH
M5Iw/y84QS5BQWWd/69xtub45SeUt2fj0uADtMf5R8cJa7QkqdE9HR6cIoNv52PUZG7ZfrBoY/I0
S0jkSOsLo/Gg1XKPx096hT5crpDIK6adgCMkbo9gh71tye1dopgmck3gojQsq66oQlJviqV/fGTl
bcPwyxXpw5st6xPW9EUkE97wQJzXymYfE+8KWdxtODp6KOJd9MRWDxW7Fk3bvPI6RC6cIdHzsJp3
rnUYMAwXPDizCq67Rk5XNgQh/L4r50vTlM0SF5sKdV6aNI8p6ckM68sjLlHQbUt1YelVeuEo5AN6
A90GZt5bmNoAp2YIs7fIVr3AjtJckvki6yzs7FWdPnL+DV3saSFfwEUvkjfc/wqCEolkuFVrqbBe
pBnouKUJkoFkhLnO/MsnwJ0lcE33y8DSm3OAgXole3Rz6G1NfzuM0m4P109l72nd6mcxCIJzpMVG
JTP1JI6Yuw3qOb9sLO+mxAlVyskN92GDykpKKh2IZ2WEX9H2zgIZm8zoGN4Vcft/u0Hb+JoTgSfd
BTrT9/uuWf81tzfRus4QIAV+OairbxHY2qQXZWj2FsV2g6M54bWzErWtJfXuaYO1rGeYVPe910Bw
RGZ5qgYeA2Mn3c8zpdn9J37leXdFkGz9NppbkgE0kfEQHHb3m6Ufh8PzdIKRWW3Y8upRhEqV1Epv
pW9kN0JQAuZkm6E2fM2p+CxpUKy+Y9NR285DXgdRdCUC42AR+JEonsVr8ZA1RGdGq/e/OPq4M+9a
Qa1O1f3EIpY4+s2i2bKztB5YCFEpTmg7M5AM3hAMAj5H+ppZcLWcfJo0gP8On89LUD7gMuwMX0qM
6NisB/KgJyWYjDHnURonSw3nj5ylfac9e/QCTsRjXqpBfIswcc1QRqyPY2lGebRKGGzfVB5GfRRH
eMgXvNHr+8qbKzlkrVrRylDAb+WolrE4VJmwm0ii4CZT2aOKEW8+XMzFBfxAIW2CMSkEsNQpyrYA
i1lEE9ZQXMstsTf2/ZSXiNG0Q4LhnzdTEuoxqVsAZ52lz/rx7lqrmxDXKOZQh2txbWzwkMf7sfm6
1gjtboH0a9ANB3S7Wf+VQGB+mDH2bwuSxJAvUDEwMQMrKRfVfPOjcL5mJJgL2veDuXyvNgSZqiMX
JyNGznlW2XbcFb5CGLbAoT4HaMrmzxBhflYNobV72T/y9BJGR2W4Q2xpcaHM9mato9e5reOx+OO0
kc4PP8NXyhimljtT75ANnTt3pgqyUmaLyjDfATa7nuJ5K56KQ1VcTtK1D32XGETwoz5smFR6xpbJ
Wm92M0B4BZdWLvAoPCUHqD1Gs+A0mir8PKDhCcaeBtpPGU/KHSi3ZHomwrKxacqfyPJEd6CcBt7x
liOXfdmSbXNp376lqpXv96G0kDrtL7nD+Wm5l3np/FzXs9xYnSs6fvATrnjZqdERCQcBdrxjFeex
DuwfKKbD5GyP+obm4QWFWoaKTPjPJrs0tBLDpzLXcmBq29wLUSbHOZ6SROu8jkZVqG6M71LSEJWc
tGNNmsMhfz/NJy8HhoxXM99lOHOENyDdCuMhyd8WEq+tgyPnmLNhCt0GSWJOEpo66p5g/3VySUhq
TJNojLKrMadZAkDjz8HTS6I7vj+3OaxUZx9oNfkA1mUp1IauYcbapKdGc5rFOrgRKrvpJcxlWGe9
XY7eQSvfF5Sph5mdBXTm5W0npFXedIj0emsyTG+/lTZXN7Z7GsUIYGsFSSDX2C6XJf/VeWiXZnVX
UUIyjliZ7k2SHEfIUGrlxrc5arXFXA9PB/UnYEkkCXcmG0pFmP/m8LInasdnOPYN1YHExWl3VSE/
AodCOBimn1l7oDH5v+N7uN8MTW6cdk4LxQouu+t6v+bK/cyZ2zTmJ23+QK4x35MP0Gj8dXRao2bR
tBslvZWokn1jTkIrgyVdilTS5hEFelEI689MQjR23w1p32Hw6kPmZHbPGhWdAyRrstXgFeJvQn5y
egL92q/NDS1uDY0AFtmhnA43X5NAwbmmRLFS6efa9cXjOel91Vk9g9kiQaZXrn8QGmy7LlWxKXQ+
ps5f0KWaiulQAozKweUcLid8dtWrhr0V0fJ/7Vh8jdwqY80gMGKrR+nIPtr8goYAJhjpnar1r/JT
FybeSvVENni6PiPOOzLcQTEcz++d8M7v+KFJ1T2CHNyTfYtYIP9gM10swC2ecowrG5ZQLZKtf7JK
tflY4K8Q1oXG0gOegpaXKoycq9gou18zwQS2eW0hk3A3b51rlRUI3I6i25n7sFMKFEuPIJq0s8G+
flytqf8m+bnjMMO/MIJ/8152ncvZOkbqDUNoWndJSV7Oe3a+z9KLxiwNegn+AaFgMdp6HJoIZeN9
uzuR0z5oSgdv4YQ+Rtr4/qBa/qeNYaNbFZEsLEP7xYAhLtqJiYxT5kiN0iytDNbViEfOKgeudWc4
PKEvQngwxbpbjlOqw3V0/dTLxWIY08R9VypliRSL+BxBnReaobv7wncQmQ7Yr3vWOkQ40ys0aEdK
FjgZjvMyxW4ewrzC+X9+fvHSV1rhzTFtw0BjOSjxs9C12OE3oIqpSu6eKlwiWpvZ4KBfJBVjGOm9
P3V5ZoS4YHZxJh4cAvG1ghNrr3LtdP9Dijcbz+S99xcUofvQQC1zgFSo5wnK8TaIIHdw64y5DyEX
VKx9eihNaz6oJf+4Fy3xA+dvQrETvlu7DRaMup0+niGkQcpWpMosRrdclJG8LudGk8UgIhKiwVuV
uMTcDucRacTKyuVxVO69NHhcZP/Ob6kxzVt0ZQOVvtKsKS3iMh4JPc4aAQEHrjHvz2muGFthvysj
zxghtDVMw8/XWiRSWmvKZj8w5qnOZ6M++IHpQKzC4s1RqdgTPRXXMxtDBLp/hnu+w1M5KcUC/CdJ
/mOuQGetskTk9ftMpWpCxevQHXytlf9cUDUJQ9PNj9gmvhs8fLKm91r+hZlbb3ZoNAgS/WmKNQd2
Qosm5zyjLqXRq56WRAkjLR824hQG4IFfNOX9R9TH3bsN3DVr3cIq2CV9NJaZqY/DlvuIEfE6Fovm
9F/XrYc+95JFAkAoR3kkOuywonAzYKWNKbZoLKRn6I6QzbflyttiIM6bV67gt2RrCswn3K7PExua
g2DzNKYEJ6/Oq8nglSwkq6zTm5B0C12pk2g7yUnCF53xQ4Ls2AoLbY+x82gs9txcF1MUW1mRh5Vv
Z8RDVt+X9IFvC0Q0/QXnPSkzgo6fry+ZFqaPSTZAI3SrR0EzAUoYUluOcSUHnGyy6+rsXjK3/8L8
MO+7X1774w0GMXvQcrK1hDHLnjLTGxj8FyEDzTG2QTzxqZZOu7EA0Nr4Sx/F12oA0Ww6ubwNlO5w
8r+3BZXoE7aOeDHEqq5iCbFU25kagGO9P5DymzQVh3/jxtG4MwARtflUJ5B7sfRmw/lf3Di/9Za2
JpHU42QhJ/OvgP7ghgVIHzSmAW+0ErEQecS5HOgky4FR8E2678eMZe0O/1mw24uPpavNbuQ5yI4x
PczqsL8P9xMQW3uov2jMTuRRVJUn8vv/6WHImEg257sqQQ2WY6s5Q57jJzBkAM+nKtmcWgkmjlPb
8qKLMVB6D6/77knh2tct8aqtZNfcGsjgL/BVe1dj5p4H6xUJITMmMNj9qxlrC2gjojVfr2gpGhGr
DH24GmMwoalhHAB3JKYzliDVwqT9YV3jeiLtQlQnYQhb3ArYV00KxGOnd2DE/FhoUVmtzYkmQ/ZT
WjHBJCzjzswf4JZcfq/lEKZTxp4B3hJZ3fWJtLJ72Wtzep/0N/Tz8igNu4RlNcAWrUr3gY4F/Lbx
OsZFGMds453bITJv2lC26NYA/seJ6pjhTPjlGgbSq8bV2wuWWzfRXdRFY7dTxULYubfyPaCQQv8z
5z31u2G4I/ClAs0CYweTWasbOgu7jcSQ7xeh9TMtHc51LrEU0WhknT+JQJW0hqqRZkPq+aD1qEKE
mivfsJzm7JHwSoS1oVIp1jY8cngu7GJdGMmJr2Dd9xTuIG0+sd4sfwjPLP0KThLw0ifH+VVMQ7UD
Ukajg9Zf9N6NSGvbGyHACd9wjPbMmx9ONAnmE98b62JpGhjsv0OcyZbr4M+UElIGQ+eOIF37eSwV
nE8mjXKk33FhGZuvTwNuHyyMEAx4sy7qWyJ2B9SjiUSWRuZUZjw5XGPYZA/8p8TfzL/TBU67YmtA
geYtjIUq0Cuuzc2WN6TGHV7oysNf8qL9bQXB84eJRKqeuIW5QZg2NG55n05U5eBY8zOeTlfVI8AK
ohaPPrlZmdJjWFYQNCpXwlECnzWUDhRAht/WzBvr3mKrER58MbplYXVSxLtMkx0g7YRV/t3xHAhm
fdyxkRFexeKynhMtCmUXCWsGBa0KHE/XnPl/r341BRFdOBRBUbPn+OsEOiodu6JMb8puehFdwZbn
bSzOg8lkvp8oxd3p/0A2hWR9AqEufI9DS5VdolvgLxJhhqURsj9THfa3PrwlV/gKciLRt7zGUeHO
Ib+sg1qtjIQSKD7N+XQTLYuWp3tZDAFI8hsRc4VhokvtxmegbmX80bImDVCCvjpPj2DT6fOjwKam
jjLuPSF9L+xjUIfWTx0CO7vxrMKQtbWCHmk9zf64RMMBn16iJoY7rXuFn0P1rHN/Vm78gxRvXeDF
FRKy5ZCbwbYKSzsplM4kNkrMnu3TyBKkL+FuDH/Dm+QCOpqPShv4h8cr5ljFf/3kb7KO0sksuvua
NAxKu4mLCzpjLUSvyxrncG03WM23osuF04Ylx2MVYFyJjiJAroI7KfCPBOZMYOx3bgfG3IEZbHGm
3uLmZewWWTV4ppwl5/0QmEkcNtnctzHVHNmUtfpeOgIzz3QZyw1qihA2xT/rxsL1/VQn3SB11WFP
kmnMvvCK+7QsZEqReSEQTuGSbWKnFwbrNyf9UuGiaY6eX+vm9iZuHINrq0Chp8moALxsG8FewbbD
sY7QSx+W+8TmWf3ao7Np2TTT1OcFu/qOlUDDRtNVQOpXlc9HU8NwllH8Y02XBDtpgIE2396eOwXP
eI9SeokK5WIqkKwbxm8QeK6o28pPgnPrW9SqYlU2ktP/uCafDlFxllXFsTxeg1Y0g2f34dAMgC4i
5fEBzaFrjgI5QGO1O28Jq90Hp6ZiKL6iEuQ4TxAuGJkUhn/8M89cBCJHpu2MHFIB8y+PvsgdCBVo
ScIgLfUVrqUa3Cu33QNv7+Y+3+gGtYtA0WbuyN9tbxwTfV/r5B1UTlMg8UdnCwcXsfuCl6fCezx2
19GKvP1VHq29QCWirCmMc7zAVtiF3pv+9OeY0p08NoUwfPQTvfoSszmbhhBAKXjefcwOHoOJqJws
vIIIUfF5XRcjzD/KATcu/tJF4WP7HojMeKSM8mT6iYISdcJWaQGlrqTVinwtnWqe7BG08q2yT7Z+
PNHs62gk0PTwydTrD3CegIu+xZ4Ja6M8Mj+BOQcyQlrmXnORd60C/OgL4aXo2zYndhdfWdFXlBtk
IV9DoeRPWzOmny5l79liRiiBfIv4lJVXZrg1Gkib2NghqtaYl5TN9Clqj67F645xWmUx/Ql4YLNk
HB0I/ySPpD+xf1+cxJDHCUravVrBgU7viN/YyYLf2tyjm9rghmvc8JXUl+8AhHXPoxvS94wD5tnU
7hYf0fag/tXnDWnW9kmxoV7Gc2rKbvvUe8QeRjLR2C8aWEYBLwFCA/izDC9YRu9u4eBpi6YZe/zN
hjW3rmeWPGgXKqiimr/iagRO6SlHLHslcIatu5ktcOjAa11sj+bdw0KLVkIY+OejRMns5scfyCMk
efJP+RYOXG9kJfb5nPAPGVYJXKU3K/4lrKCqUiOFm+RBDxH8Sdk2546n0ZxH6bj0jpjIJxhR2nv3
dw3QRfMvXlQwYjs7hr9Q13jTZ7vKXxrr7/NyZKLwyWrDIZafv/P0pHZWecul81Rx05zRRDdLqdB5
oTK75CAlVK5mN0sP90txbHDpFr1KhtmUyqKlZwv70DkCHePx4kRurdxj8oSNUoSyNBDgMoMef3qY
Z23ryL29ZbD1ULW1/ni8G053T0BVK/9dz8+En8q5nwdUjuYl53WFrK5nYrVFwCtuL4S+vhNT8cG4
0ybv0p9sL98HE4BTIa3wbVJqpvMEOauVJ9mRrOPaC8UuvORdbY7H+JtEFUSJptFtGoukuww71Q+/
TPq/oS1Je3E1/N8YmoqxuOH/hEwIzdfCNF9XvUtppZ1lsLGC+ghsp1kM5ghaZfWIuV8LwKePhBMS
oXxhLhGm2lqu5JsbRM/JS3GqiC89+pp3hI4PY5ORHmj7quhPZTWB89s3brG4/DQ9rrbdDzV49aJA
d4mCiqleYDIJRWNRTFJH3C443N+iDHpES4AgQu3Yc6e2ZRRQ7uM1KEUxhQzSyCZWeRcc5qEf5eiq
jTq65ap39UB/GYDxyKfeL6o2i366XXes8O83GsdCaEK5eCaWKvkTptrk8eAVlUQUmOMZ01LLAUuQ
4WgX14/x/7DmBOshumkMDPd7KWpP6SpIzSzYr4lTILGdVAazVZ7uUbU6OpgkSgT2Qy2/7VT7W+Uc
Hdd+tJWASnzGbBN9oBU2OQDyfse792gUeWr0Rqk5NP+FLRUm1rqDhi/wTK7q6/bBa/6SbY0mmuUv
A8rh7AS2uHeeVNA6ACzdumsgM1ZAUZB6T4djXRRdmTCtPLKjFpocC7NDkIKNQWuKlDusCxpXQoGk
p/LCaruwPwpVbJQTFp9DMogx2sKtljPTDEcfsJlY7LrPG6VLv2g8sNfcls2030TD2f3Zmr+IBLhS
31hY5Io5gWny6xXLq7KLVYULGg8H2bKrlP4NWLE/ZWPYojiw6tZnaOTpszvjlGM+Fk4w/0TLOVtp
pi3XKAm1ZHhixocYBRVCifRI+sRonoyouktzip4bBf3+CDZ/lE/gpL0nR04X4aPGUePIsgD9Zcx1
YvPv6ZIrd9Vh8mRdAOaPV/SpAq5KkIUMQB1BrzA+iDr6Bc7JbIe/9SnM5uIDTm+iF6N84itiA6Jf
AmnMgiWvyFA9dOxopYKo0J9QnHnz/wriGFgrtaw1Z89ATEfq0coHkJQHC1zrLLpy9IB/N7zgGAku
qsg3/EAQbAsB6UUv0UR+4ROCNEuSSuq2bTFaa52GeS4uKOxllzTfqPlKbGxGj7DZcl6RHIEOGfb5
dqbwZmx7qZqtA7udQQ4tGGf9YGggseiUm/xaLGVGNqgLi10xH1e96n62Oq7kA6VoKUIaRFgsOP+X
bnmlRHNyZeP97IcCCjg265W0jSf0gJNqDn4VyeVKyl0Aw79BqtBhA32iHa0NE+nNYo4/NIlaQRvC
At8EOul7zNWKqGgVazAZ1oEVuqGE6PIDL2tW7X37aBCcEFXJtLkQAqmtgMWogz9zYKX6vCdrl2yG
rEgIGV/fIlmGyFdrhoc4gVPukzVC1BZBC95JI9yvttn7gH91Eh3w5ixt5ZeuMWE0A+v+ZnOjA8ho
hq1GjNf4gQPQ4uhLdEFeEGM/ZG95HEWo3mQLLgB8dD7enpaeGoHDo/C0KMlp+p4LOqKhFXY3HS5w
SlzUsosGMQURVMH04hDbmyg3Kj4hnM6jUTxNzIl2pGeMJuntvfnmsuuU08H4z4PNTx1tpKO4pLoU
6beizs3O7KD/7ShVfvahphPQySPaZYiTRhZd4idVwv/7e63cK0aILt0K7IQyB4c1kCserR0yK4ch
wPzxaziO+6IVXwQZpRJYUchtUdbs5FXUYEn+PER3qo9F+ZEBb8hA20Wmfie51L2s6KGg/DTQHjSB
Ous1EsFI0gq0mcbtBK4Ot4DAC92X8FqkAFMSwjgDQi7D7ksRoVqyXcs2gMnN//xABud3U+7u4zyc
3RbNyZzxRRUZ2cW6zJ/2aOjUPal/CsLZ5UH4+CmswAf5AzATETk+DSzBTIPsoXH/VnOW02gnWatg
7Kg/ZphotDVtMin+qgZnVMOyxcFxbqsz5XTMli/gtA5bsfItSVIMyb9H0YA2Qq8yUJtpTpCD060z
/5KGUuWGF2gL2LoE4bWyNJupy7p9wyJfMa083j211MT3eG3doDjZCLM7xOYe1Bde1vEOoXxOJvPz
g5pUqdrc+yij+G9jmd2PMZihZ1N0N6NVnqfzYogwBAZKcdSt/qstpvkiDkZd0hL60bW7Ps1+/ZNr
CC3eVs43azUduVaZJ9r9xx6ulk2G3i8ix0EibfMDLgNMK7HuTnUrV5wtuGu4almWFHevNIsaLAF7
jECiZ7iZTHSp0OXHAa3yPQyP2wHzCksr4YUMV6Q7lUJ1ich9dD0QEmG8m9HWpzz9nDl2/J5+VLz6
Kq0O3wHmDOtITRcTBI4XCuQ3aleFql2KbocOboZbLi20kCU2g8XTI6dor0w/B74oWMUzczn492NI
ereA2SnMcjROkfC6qIJdlpYDFq0NwVJvkZHYTgM6ZrdJeaDhFsRwseX+QZiQz8LTSM6BSIVLuYXn
UZOzjr9AsnYyWNL8q87D+Ox5LFecRYYK7QXMqz5EhTUSgF0qeXxYOMs3k+ydDzJ9pItV6wjoiBMP
z648/e30JgTVDd14gjfLjLQrGV5CE/rB7snDS1jD3jbwbAOhjLaW96/83nJOhMrVBX09w8quEZKX
sJJa/UawaXeY77WuoIGnWv3o8S7PhjyBzQ9zbXkhudOPZbBpx8XcIwW9lh0ASxhMm8lYrEFfrreA
ZT/g76+Rq8rljyAS2cHrrqdKnWFe8sIMt1FWU0eug8Gf7XZ9ryDdQaP8qwZe4ue/yD55FWJJ3nnV
3hBQiZnBUcX6tD7sHSx9fQvrIyT1/Not45aaQd+xomVkDXlEJJmH8FKFEOzKVtnz6zSuskbXFcrD
kMVbRO3oBThJZRMqwYa/aLJqt/SdWseJh8XpyHof8Qh7JJCm7VVBlBD7O5DF9g5E7J3HACWEfYBc
qXcQLwU1dNFUShUKBwuEQp/E08dmO/5EQ7i3jJH9NvH3D2M8r3sdWPckccM3VHQxI87Q+n7Nq2s9
qOun9DGBrzoJ1lmi2RH6c0TD3mOVx7SxKkRDv7aJ++rA8ZoOXBGTvLF/yAybKzgnMjXvmp+QDkZh
3MZXBt6UMcKTyQe5PhtwR+o26IGzap+3hVgSSHgjav69LeIzlh2nOfTlkvO+PYDppuDMDyZ9j031
MVEMG2CQcQOVv4cedn2RsvpGIUHIxuBgMXaBoFhrej7LkvVPyxuvJ+2PXs1f7az9oMY/fnJexX8/
+Z2hyOKymXrFjS8wr0KO55xFc6cflwHLc+4GgHsAo79qfJIPgAUmFvqkFf7gI6GP3+vYAyOrYp50
IJTX7j5bYexU/y2aptbolZzPdzxt81YntYHtbdTodDKDANkS+iEJ/cfMGZwyjeG8r3TvykOPUjCt
rWmhiaXWVJ0TI1Qt7dRvJb/lTrNY3r5GcVr4yWo03wbs40eHIPT2Co1iYjulMBFylQwfBxnVeCOn
PXKsmqPGojO4GRmnxj1126qXzQsYnJRyCqwdqoGSODMi67hEqyhLmnDfJWuKYSmVwJWw2X3b3cuc
mB6877WAqn+KmKDRY7Wp57CFf9TSpE/X5GjZ1JE17fdyyn0yfQFtrIkmMv+5tW1eZpbhCfRCUVVn
EqAGhSnWxBuDdfyOFXsYTvN+fczkhFcvaybcTJQ18SkBRNLUNztBd5uXNAO7quG/aFLQgWs0LNdP
crNl41I1NitVEpZhZopFXyuJuuCC/1MBOL+12Wzc8/0Fsw7QMTaBZLaE9mXZ28SaFKn/8P5L5n4e
8mCkmXFuF6gIr9oxXsKkrwt4YagoWXQKqvdrxrKGsXP11KIKOxc1sjav8ZB5LS70lTfcPljBxgbX
mK6Iyry+xlOSL7TcGSrfQhGmeZ6FY8zAWhWaV/ULXzvwqjj8bFl1hMkZpOjnmRZri/sdX9o1buVC
2ae4mCwSP/ue5wyFjQE2vph/1TpJwW5CKch61RnEXCBYGu6nu/MDiNBAvyJ6r8bid/v9tauM0iqM
0LX1TBtTkMbRzbFDH9Jy4EoLpKj/nboARD0Yu/0+Qm1e59gxhSAS1vnTpbjbUXAFSsn/qqr1ddSt
fO62Y05G/MFwXRd+Tc/DLpk/ldYuUyZrVnpYaKt91qoRFgpfI8W/SToEtUrlhFmgg+WdgVhcqPfO
0f2X8NqDcoCf6E1xvd4Q0uGjLRuvXar30fDLeQ+Zo1xIgPRk+rBuIYdBITBUnsq/OlacJCp6bwFN
tA1n38sq5Gu0wmIXS4nCykD3EYOqSR/Op4u6ZShiDnJtakne5/dN8p6kkFx82TpWY85jUHoiOvex
bk5H9VVW7D1bwu/RZ1SR430xRppaz6ludDizHn6oVHzHEhcDQmuJZ0P2soBZXPgLUcHG+lxad6B3
HmeLoZFrBFynALGwI8TIhUt7iI8bgGHlcJBB37sweyk06yrgm8gaiXbvsIRvRQDhfgs4PbrPs216
NMXNfjVc0k3C2p4P6vL+sbKF/qQaQbjTvfaTwUvZL2QV23bZyKpfoHllLsDy5VbeGZQ5IHRut8xm
CzH7LSm1VvtTyhD+gruO9S1YbX4ZoOExA6xWyAkY/zObri6q5VrgpuE6CuTUznLZyZoikMWF3fQi
1Gn9VvQwDuqJHl+1gz5QhO2bwqCqBKAaR2ov94uFjiWT1WirSvWBRT0zzJBl2w3/fF35lFhuIYfF
7uhFLFzyELbbdgnXlI0KuSiFKZvVRRUWujmfCQfH98OJ6Mk8wCKnNq0EEyfp8ht0SlTg6SkYMuht
aXzfTdc4dYFaOkkR8iEvtp1QIx7PnFz8kPd+EGooJpeNA/aW+RT9MdQ9hdKkbX5LqEu4nQINLDl4
H85mM/nPTDYibhhVLxUh2nh9P+v65lcnRiZ9AGq6Wlr6T6IlF9gw4fr9ikMefxFUMfp1VoGoBEON
F2DR6fcaleSuoaXVr3VThJpHc5PryqxMRxpepuaDLzFZy1gvMIr0ysGcVqRsL3s+Yes9Xc2m+P39
iVhImfKqbxha+n7IvcBaFvgUd65H9/U2prLdRvGzTA/6Xvtlm/U4xdSDnEl7gjgqP2flpqLt+V6g
bTokwPU4ngo9jYu1tA1JHiSmazGHjIoK5I3UB0O/Nw03K+jBfKSfdHcyhgv0DuurmLDcgAdAyoTA
SsWjb+Ax/zPVlHG7e6j797OCqrIkXn3RtJTov3fiAaQIoKHNEpdNcaIsdCwvK13kMIL6DV/8euuD
G8iC0iXySGhUxiAGAxLtPcIUoNp3qVqZe7kq73YfQLkl17b14D1JwpelCuc3j5CIr52T5QCfLXC7
1lGgbw2r0ImUMmQ5ZW0lRng15lsVA3h6BAz99BqZaD8bat/kPRiXLq7PAynE5NGcxNvvEHFKoCUa
MK1LKxABilBpi2PWbbQ/8IpclGeZwZi+D704hIDomeM3KPfCkhLsHvPWfOe9mL9RQ+KrSt0ZrBoW
gOYRmkiYGAQpeJasuqwQqevSbWBVY5KCoAUgnNi0+YQb8wXd1ftdqB4euwUR7lLf0rxiBg7WBo6N
Oehk91EnT6AMPF76UzcUr4Ovjg8fWNft9xLr9xCKKebXeBf7XoxwVFjWW8djB+F4XbAt9ackpshF
MTtrWFzxZbeddyXN1G6wZKyZtyioBsGDLIqxOWQ4Bawk4hyDLEeR0Et3GVa2x8JqYLfqUOZlASQY
hJxaiX8bV0RO8iNE7EDqfaeHtjPQal58IXrtkrrlijfNZtZfA26Xt3u7kVUR3tqhOa5Xmqm5UFcO
gRYeYNHxpQIveYGPFrDpt7IMLGtrjfuQlAuEvGMiGCkpBYVHDgO0RQrXWDfcc/LK8d6gJa6yAYl2
zlkLmWp9NivDYp15iwTtdHkutYVg7pV7hntqj4tEJLnd402k4cNALWGDgzoFOeMkfX21G3o6wqGM
5Bz6uH8rO5EkByHI1TKMFqv1jC1FRAyjpmqKbfehXJKTKKDgNpRx0eRW7SgSpR98YrA/on7KvnLa
0WESLSXQwoTv8bgY9OtP6LwJPCEqju5yBPu9IB8hB2CJ6iJrl1XH/D0ss+1QN0zmMA2soy8VNOAW
vFxY2um8e7ixQcM0ihasvAt7kTifo+BKMgF9/TogU5O6IsEQl1DvcGN3Dx8tcr68wXg42EQO+afM
HCvHxfN4TPiOeecE0xQBUOFthN6ED44wmr2WfabnQLBVX6CPKb2w11KEDoPG+7m23dfoBlqReb6S
j94P3PTKx4amX1E7W8vYl/J+TDFDWZbijD9inca2JmXW0MNWKnkVfcvMYHnzUnb2fZRb5wSpNm2q
T2ZtEUOGDNSDyFUNRH+C5NEydPPZbRdr4HqvPFUsuqVKdsmXTCsdzjXyX8jOrY3MPlG/+RPguubJ
+dZ3OvIZWWUd35ff+1o6Io3ULMVwvXCnbZyH6N7Uu6N4aA0NW0lAPXiTFrZ9FXaJqyuHjdpg/XfT
PXxr2Xb5CQqsEN9eb5LEcHfSdPtmjd6KVimVcaGwTE3WPGmtATrFbcJhUK8JJ9jYvw6jPlg0JhkZ
xHHuhtKI6k4RFg6QoTogzDvHDfxq42PO9S10XG75i+ng5EKdQd34/LUSzJq/Zte8CofDKvtAs6tb
6pktm1elAblqnJisEzH5pAaWK9uTzSipK5sDWQ2DLWNjgvCKKgJI3apk3hpxioU4JTXirsXfXGNr
UQ5ZSfY5+T4OMcZyZWx0lUcxCkEbMzOCb7Hs7R0cqeQyFXsorMcZhYJ7YpeBovcVhOlH+0KdwQ9f
jE69R+PLIzd7rv8ql+AxY5x5h1NCHG4h5b5vLKpupCHbGvsJTQUGYe9K+ntThiZaKhrZFzFq6INt
rMXL3rRxN9xUq2HFQ2FKcrROfbkzWzid5lm2dWtINrIH5S8YGrxxz1vHWsRpqJgoUHXkgj6sfZ2K
k5VbdkcRjMVzqPaDJkA0EQ244iCp7XV1AyRsjA7fxgOIqHyKcdZnWeTRuIvKeuwQRapgD18r13/u
9GWjnG6N0He4D4DPyuPtCSmtzDkz/Z+rf0WbmUe0BNAihdjkmeB0grFxkiQDQttHxbxfu/iZhulS
AABuX9bhVMmNmBwe08L/R/BBazIDyHpszMA2rfMeZqbNEb8/8HQ075hxi2oPEUGDIp7sHnewihRa
DMy5eDzPhD4Ra0fM3/Q0eeh5oqI6IVaz6ZU7tLv4Lb2T+k9wNk+BaZE2G6f02ARx1gfu2yMaPYb2
MRAJOgtCwg7m5Y8SxVz8W6NVvGmz62xyxbNjZfKxij8o+/p/cjdg3gd0UEmRwK5X4YfNo9oo5xS6
48EyScPYXfz8efMbUPOlpEtoMEEdlA75fZV2QMlYTTUgkQHMJlq99LAkRFoSdZwQ2nMCtz4JxRsp
CVx4iPtMpSZP7Q5x1q7PKqpa+O06d+2pKChfS9DVNjF2XNB0BJV5dUAB2pQXwEjDVcsvJ/f46lDd
JbzdEfEfm6S39M3LaNGwR/8MBZNUzRMU3yiVEHeyce/TN7ea7ykYaZ3iahIHnBbovJTd/WpU/AZO
5u2ERX70jTRGRvKcwqV4GuPa+0uIUWL877jskZpu94i8ftjT13l9RlfMXU4t++R+LzBuRT0EBJS0
O1NYVJ03hhcpcXRaNl1yWsPaNQiv7V9suZKyf/fvakV2o840Rid7Sv4pKTiRUC3LexVT8pKSbdgO
u8CrzdPoJZicveY3lA1SDHShigflcHteqwmklcN0xHoJVue+UcKmV/qixzeeVfnNwRBz7SOBt8ED
pFCARITrRTmMHANyB1Yx3GodaR0qdplCEVfCc23mx5yKN0eKIv+yM9sZOBfCYQhFu3qDamNeBxA+
PIjoUB8RCEW4BoSFHbxuHIJgGmXPNFHjcA9v2JoZ25LKlr46ScJgBQe7RmVICVKhQgUfqJDEXG0A
R6CQAzW+hFFvfZv4HYhOFIdqABjX+9w+YSjfXkXpfELo4HrOwzyxEvduulk/V5Rg7iJW+sVDHijY
sCbxSJeNUc2IQeZBshoZAZFCdfIcbzNysbLPYerm26ONkAuHANPnLUNJEPk5kN9Ne1m/XYJALwgG
1bzgQXIqxnikQpb/CthMad/l8hDG2U/9BsZLmUhZn6fSJf9+Dj7fixhgTz9cG8jTlNnZPg/4VflW
gUaTkJpMlHNLElHhSiMllBHH2Zw/zXza2T6ZO9hS1eDyKjAKGjgjimjRwZ7472Eug1+M4zUd2Hry
kPMz3wfCXt04JY09d3kqsXxHYLAuXNVDzxRUV8/1OJEMrx2IJ4ywwik43FX6AfB6oAo2LeNq30k8
wFzmsTPKO4tLhtZIorBae1r6JG957zK1ZAJzpOIpAmo94HA4MrT7xaqkgXOjzakUfdw6TPDoCIpC
IpUuxU0FGM2Cq5P31UwiEO8HAIsYgyb7Ubaws2pyHbNWxJxTtI1nidH0PLC61V21hxy7obMICO/N
xKdr3y7P8FAq+OSebKqLocUpN5lcc6Nx/gThJJM0WXRjeIq5WwsIJ0aRUfhTtw+rsLi6OLun9XMy
hQAVoY3vPPF0ePKbD1muytsTs8Q3cz/kXy1hZQSm+lhYaDdZ+b2GrhQLsNAQpXtoJXjQ9tEgDvum
6YqSJahwEXb487d4AI8rgXzr1PVI6rw/SdZbpwDmxxrMKxVyY0WZnNr1ZzxKKrlBxzjISIWLf8S/
9d4e0oZq66zSTVO6YOSSIEzDp5AlBFQi/R+8T+LCR37A1ly9sG4nZVWgYgIUBKSbv0ZolrxJkDFf
bn2ubrGZrOHp+Awy80EezZVGeaQk0mOl0qyB2gLlQohc+QsFejdTCqS4SXQtYJf9yMmu1RUCTDUm
jcS3LSz7n7JWV4Fq6aCN1uvOP3e+ym1wTxwkxGYDi+rAMtzqaPYziFJA9/eyYrK8ODUlNtKeyZyY
cafUN8YSeuvqWSLfbhRNHos05q2jUWLjO/7O/t7lCs1bu2pUWEIM6khmC9XBdJ7rrM9DUUTe5aQn
ir9VSgVmk6GCeMl8g11XxdzSX+diM4wRJknO4yN0YAzJR4s2ejGkXaDuIdg5bmt8W1T2w1MYPlQj
hB0ffKIRSz+t2uZKkbVR0OBwv7v9xld6q3ep/8ekfjBQKu4lRK+/DIAte5llyeTFx6KxvXr7W0Xd
2mIxTOEaVlzzMHNsBP5yIFyy4f4zbTnWd3nUa5+XovEMhsEYl4+mi/XQReebd0t7RyDKZcaXwKj6
lN9Pkxr7Wx8Vsx0hd+e8ruNeCzj8I9Gmw2T3CQxQ0tpHDTqNHukefUW3+kgz4vkMFgo3BenhmVq4
LXkgN5G9PTdlXCf4rtaDACORuRUN3bjyQa1dYEeRL0qfJgHahCCziX4XSX7prdIPOcF6R1KHCABO
faSM+LjqbVfN7iStnf+Oc5x7v59bRFjw7GgBudS7TTpM8cwKSOwXCoc8+ai11FhDgLRebkbNP9zo
CpWreN9lJOVxh+wy+iJeKX6XHr+S1dJc1i5YGxIgOA/vluCxF1ml+o5Th5KG+sO87u9p7B6iiOJM
IPViQ/CkiyJKnV/RZdDP3SIzOqcSutOSyJPxHqJdjYrMZJ02pDSmb8cwA3A91QFS/RujzWyF9jfb
ly8hSyr+nkDwcZJOmedfVpLu3hKDJB1rzMcuzGFcnVaC4/5rgtWqSLetTwhRvHX8rQLcBwIm0Y2Y
kMlLXtkgkGeHAgA1nWy+DeGbai2MzTyxQK+/u/gqiK07OiSHAeUG0DLxT7J/wWIBFQt16MQ1bSzx
5TCb6MCIN6TFSsebeX9Mop0GY+kv/L2ZVdX5TLSTxELPlsYcIOwrZbrYJ0h3Yvq8Fc195jqVOJkT
orD2XYIq0rDynCkEG3wsTFKGPaBCujfeeIncJCcfJPhsAAwnqy04+iQ+EDtAo88LZs/cAijYl80K
6yUaWBNF2OgmbpxvhVivpn+c+xZq8G2FU13/NzHlMXDe9t11InpO82vnZcnHcqY2/St/Pz+nS2Ml
0LreHn7YU3qpjuN7Gp+gJpGBk+SNjy0JuEPXYxLPVsdcBmaqmq2UcMc9KQ7WH5+1iDqHJ4rNTd5j
b1lpDaTPqcahf7LiVkq7pgj56WPTQlbCHRQDxPu6IjCGRwX/aNP46bNghpCFcPk4x1C57HBv7Tfi
MEtDHg0LrYVZn33dVzDHor/Q9+7y38BxvJ4tC65ot290wNfunEJ6LvFBZbJ2hioDAo+YJAPF2p8L
HSNhmgCom/7z/sj/kk7Ifh1pF2jsWstUa5b60csf1kgAid1SpFsSM+GJpYRG+9wtQP6qi6f4qrOp
oxbhVNA3LWuSokLnyToANVhBzivYK2heB2203f5ZQXFGAToG4dFatQaCjRZz6AS8nXE71+/j7nGJ
qP9ntTmb6oBu6tAl7fqTFhv0B3pQdipZlJPfHC7cl4I/4Nt2ru0eLAzUbkVZdmfQvIzb0CZDtQ6Y
ESECyI7bL7mHTlSY6IuwnetldvGYjK1M02GK3CLvmhxZBrxme3eyHZeM5QVWxpHunz6o+b3K6LTw
NzXETttv4FVbFaKDYSJJBmE07f2MDcAV+v7S8KM5gtvXz/vR9L/617AlUbfEJwAS0GzJ09nsYJHy
wylaIwI4gKi5rHsL1f8OIDUVwlWwg/rkKvwFWlnAK6rVs4cR16084ezscHUjuYKGSw6IX6X5+2IK
ItcvlTCN/1lIXlpaYNYfzHCO+4UraQF/9a+v9bKf8QYB1TRGM+qnvhDQ54Uw9lvdahYb0mtclS8+
7udEa2Du2XH4UQsaJeyAv+vQnawmip8Owu+Wv0b3kvx3+b/oCSNxTZPBcsHcxon/oYlbYYPrSr8l
BlEkmPgMHaTZWS0tbGjygmF1nzTA9nOZLr4Zb37M6uJQNSQp3jeo5kCzN61DJXEcM+fMEkh/zBmB
+hCsBZ7hKjb0AHUzygx6ZwkeoytdMYJM2ljXeIYxXrFm/kLYWw5vxIW21AgsHbo+zKRxa7CBYyI7
W0HnXuVQUwN7QU3Dl7p5yhD/+ikTtEUnvZrzQR8chr1clJ0LJBZecxgCxHiRHh6lBs9x5N48xMCx
gNFgg9K00PBG7TZcwSrSvkfagKu5Bn7+POQx4JJr9t2Cs18q775ZdSf7cAXXkmdMjOy+93g6PwjK
/RkkpSYxEs8V6iIvHF5ZBzFlnHNoJjx8TtNfRZH/jInRZ/T8YIzYQoK91wCH/uGzlVFqNh1UXuXx
torQ0dg+OfT9LHnS2E3J8/CiADD6RbwW6zNjJOqC27q+eVfGmwDRuvmnGma2Btv2RgRy7MkQHCnr
hpyQWWRYrS99QoiVHisR8FvrqK7JjX6N8kYUDQe2V7haK3RavIis0m8mdzJstchRyvB95H2bQFAr
At0HxxWaIXBD7l2mslnjmdBknHZjolZHrcM1VqmLBHmEo3hwKoZWibqPgirNWH/U7oCoC5SLh2uK
Z9q+8Yl+v8DfCEAoHgbIW+WYiTAP0/uZzG3rRf3TN+BZcBFPfnTcpCKK6EAWCGVRY0bMnHLFd19o
4bRRfrnfflsu6yO25KU6qBt6hLnF9eWX4n9j9ZftPFk4tU/5G0X6ICZEO4Cgh9XxdtJ5kqSjQ08F
7bfPQI6hIzpgLREvtMgWXBFBFy8/jHx1BqzG7bcjCS3debb/Jd4vpl2DdGmLaxn54pxHsmT3B5Aj
mxDx1uVmMLbBKwyVBwuzrKeUEf9xEJNIbnuXbIys8FQRpqwT6EPnmfa8QqlgeaN+vAJi4RYBeHlD
zNTTmpKpFklBsICI+lSmbkvi9hGcAPwo/1iBfuavjLbn+Mh7bbUyqz0KAKSs3TKLrJBPtoHIhRHa
cajogmYxqoD44nkbgfBqc+TiLLaFw3KasIHOpoLHdfYiGcKGWZBCu1d1kV5DDqHfY5g9Ai2FS47O
iRjxeodel4/RPnj/N7UCSUQ8rLc75wc2JUE66Yc2qdYXnCrhzo+xWSPARNTwICEc+H+RAmYGO/mS
cJLQ5NR9dFFB5bXghSwFrN7u6tyALU1cLTIYMFCj1QE6pw1gFuXGOdcypzSLJTUaJENzZuqTrjyd
4wNdUv0T++H2eYqR2O7hS4HtOd0Hg3ZFeiua/GOTDk3QSccimQ9AWqpKzSHCNCxUAhxqDBUJttD2
vnGAS6vICgjhxekOBgzkIg8au2eF8psntRvSXnmQtdzg0yfOKKZ5h57SVbfP6TSzFi4bz8rc2S4m
MEn2e46IFmW1P3MZs+OWcH65RjxbHTuIHjJrSJBh0i7Y9xL5hPUFNEhh5cobJaPQAuDYYDE+C683
6j4CbYmPO4b9IXaiey51o0slpCdLYukPXMpE2w1ZrLXLU/CMgpVfzj+9aIhhXXsbWLIA0uT9nim2
O5lP2h2yPhfz3G6jzoyJ94wEVZbW/RrxIA4/m/OOx1Ynbn7df16e9i2Pg3SgGLv/kd4K+Z67eFJH
nlOR0DijJdgJy9Gpqwvg4TOzhGyp8rtxe7FP/hL9BkJtm2xUe3QJT33FDmlo9t9vwUXyCWK04rnP
CR8DTLo45XMr0oNIo7JrqZkiiXiD5jG9P2GBLQtbYIQUrh8OK1weqF+soKDF+3USfD0L+na/34oU
5P7badXO1qiDWOqXx2VZrNe7Y7gKEMl66I6QEbyrsSTn96H0xmTg5/2dhrdd+U1+fppxIchB5Vba
4ZMNVbQZSt31Fj+ZOsarwPGPboMowVEqPVEAzpRS0gXX+wxEhy0Bb4X6FbgcuBPxC3DHa+c4V6Ia
3RheBFRdGJt/sGaxOPnwBDeObiu0GDLOl5YgraojwnTg7+ffi6x//cI+aom5r8dEFc2dlUVZ+Axd
1jNkykYTddI0x2jA90/wvQih06G4BiVeW872B5zOlEFwh43BJtWlKA6wQQecozuo2d8zFTe0J/MV
F6GXrnJW+oD/WphcDGJYB1BPUnKmAs2Mmiuol7uJQ6MGVzpULt0wEMNwG773HiaEs4n62MWLLHX5
2dZuglsGZwK5oIKs3cDMdGcm+gFNuDCVzlKENnNccMYdY9I2+B4xn4BlI+4d2enFTqOIpVnyZawR
t4Ps2e5j82YpxJVeDdXEF7axr8/luVLc+rh4dMm1m0gQJiwniZYC/5TDq3aARuzxnUTUexk3/nD0
k3Ja36owtFkJvQnMI6+Kq/WCEPq3TEb47GOB6Oaw+fG0wC/0+HEfYKMldkxgD++dFUugLBbkPx4y
/1N8KH2wr7zw1QWdzFaw2xUDF1Rqhl9pyIxnilLSs07Lk0SYjwUwPskR4mPRbre/4z2dF+di6UT9
+EsPH3KxuUW8g5QMcKkgfZXqnaIBbjqnTm6jp858nzVXVSvSOLDLeUsd4NhIKLlYbOnnVCp3d25i
pfsesDb+yJlA3zY99O8JaZ9v4h1fBCxd0VTTxX4F7RqC06MwxoVqYVfZwSmyt9NKqAmzKvJ27S/3
rTUK3O+oI23Iid+lyFuwcK16WjTp+ByfJVhjumGQkPC9CQD1pkI3WHDyeoJ0p31KXL6SafHjjdTD
jUCTyl3nhhnYrgwH7A1cRgyN5maXU4NevZ6Fe5IOG4xyuNScjaMf/QOO6WB3Bln3xGGcAhDytQ9R
FcN3f/+YKJHS8Y5dLaMeqQG3AgpXoPfUgxuN145R7jEmCcVK/s96Ray5gcJnvkoMqIfy92qoHpVM
fleqYx0Ucn/kivlqegJkTKbrNsM62b56Tnabkkd+4ntaVjaMzzLu82xDqNfVoFpo7giekPk2sFu2
s440qGOC9tIy1OOL0D865rkEN62HkBOndOVIM9ZY3ShOpgr3YKAZ1S7AMzWxI/PUgLKUWuzPloJk
j9wC7f9k5q/hG5m8DKfE8Q7UlHLvu8FX6Aceqe01zQil5fHpbGC7Rd3W4I+LPEoCU7dj3ISN/NGq
H9v40gqnIvvnUd2irGDZDBGoxgFQZG1dr0GuwWo1sAkxvjLtmwNdLR0Nt5+o76PNzaqSJ0NCLvXg
/gFQ3/udFBWSikRt/8EdLEQpQTTNVPlitIb2VSBs6lQoVk3M6gljr4/KJ8YRlMHWVa+8hYfMPfaD
oNZ7UV+kzvBO3yy3TH/Ez8gskcy1aTxcjU0gLuL5lHHgaY3UhKO6mfl25y3ZdvYD6zhVD4iD3Ckr
vZHv2wGE9G6sFVTc76ha0E2VYjyPiO/1xekqOSkxJpgmg7fIEQJeR/XO9l2t6Q/q7PNT+51drNRZ
5pfyH7w0D8dKxsqf7pfbRpRkdfOGUpw23uLu4+2hIQpJsNiNAhESOK5Sij00f++kt4mRTho7KNxL
H0YqjpNP2/NjJJN9CfNYF5Gx8KB9wd/gctF5YWASdtr6Bvzf+efiF5shN59pdhMdYq3TrzRGnQzr
B6weBLjcFe7ALxISGLmK1+hBdfGfWgT49D1xoHHktVwAqTI8MdN6R5jo93knlUYaMNecUHQlYkoi
n4FniFYmCP0uoY1ibH81FfjwkS2ddhuRWycWRp1kkx20zhrsWgKV7MQILaYyVV8hRlKOy2OZgsa0
vtqe7BZ7AiNpQEwwHzIjfTydH1oCalFZAEczW1TSnppc7mK9npIOd7d0uLpMRqMfjBOmFMAFIUC4
IEumjRWqM51YKTcy1PEU1pIhgYBnnmf14H5kI7wh370i4eJ8AIvL4FFCreWfjxnitE03ObKuI2xt
pLyaBn56fUySJINnwY445+pH/Lk6AKefhVxKjXCu6HEjQnZrlNohxQTaJn8zfhcCSJfIJ0ZdgXTi
QLbhZ1yIxGu42rQX/C8ZTY9ThgRpI2HDS2XveZnzkyksJa1bVTaxXOh4uDTxUX4YvURpCQ6REWTL
ulPp2b6d6/7Ywxl/sqcghTvKnpyRRpRHuo02QWjtlAoU+M2z7KrwVkpMXiEBmU0fy8J19OwO4Ls4
8Eb3SHUAnxeHH0kRBQLyZjnxJT02ql9U1d81On5hetFic4T7prftaSIrOrP9NUfBFHL+O2gngiNK
fudMbwLnEYSpU3FJCuTDSaHsFUYg6qJFx2Y5j7fJOpqNsDnxdTO3w1zWNaOPMVLLULJWY1+y7/n0
AGQT6ogNGZ8n5ILI3Its4cTmfqnD698YL1N4Zo381biFDmvpi/YEikrqlHX2UxgIzag/hvC3xtjx
bv/GSCLxynETO1WkCKtJ1j0RTGlxNzjm4/MeO5e59w6YiqH454mR7jOAP63MvshGugeSHX4ikTUs
qUmz9qYuYDAMt/1eB3Tuq8s3UsjuCuy+ik1kRJXnqA3GYjVzzTzrmJnJzHsNohwhQDvYGfEC+MPt
28ItuQktibpUCJaw5a1Fd7C78y67LSrww+OwFBrpejuxTqDXsFrKjM6J5k18ft2VZ3IJCXn2A3Ry
7Gg/IxudgSGR1XxhblWi85OCrGU3gm8mckNsQKvFsBVyHJsdKJx5Pw0S6aTSvkMoe7cNNkYt9Wdx
OZSgLPxSVnX1ZKMxIXV7JTONVGgEuYIj6BuVxNQJqICx4SdwdHuBflbbV9nX1ZC60pMIJfNY52HB
gdlPvwSU0rtD7IVmoMi1YexohFINSU3eQAmhbUZ3l6W7QU7MOvipz6nSqjp1Uxweyde88vzaE9O6
fihxjZSlNuUW6dMcCoGRQ5ypWcmVlw/lcYWdTkM2A5utC5A5Xi6FKX8alsbnjm6Q2TmDtaloVqdt
Qkg+BZLlkXq3oc/Bz/WmncVHQMbgTCiYqkwfHnoUkGwpZa1ePN9LaH7pJukqTjQkBel3EyFo/Ytt
CltoPeBW3XrmzW9ze96GyLrtgkfNaa7wN5DxjM+nJPnexKRti13LK5bPe+k5aDc8ECgysBvc0g3L
Cr+khAWJF3hhSgQTecJYLnrmpTea/3avLOeyB7Kp7k/XF1It0e04DLVjbXCbPdEy+IYFexdcYehQ
DA1M+EqL0Cio38uHmrHGC8Orysdh+ugG/La2hjpil7HoG0MQMeph+FvBWy5DF4EmcS8eLrntK/rY
/7UIx6nXMcBVNeGVFVsqAsZR9XgdjgXbh1g0AfZDmCBpcvNqKtu/x/gT+AcYQQA7lKYGK7F8W2dR
WDQVworjwO4njkeeAV4QSrSOsJsT2zpvCnMiIilOis+3T0J873pA1faofPsXKdNdotS5tRJY0SL1
BPhQUAXaAd/AcpX3rttQBzLUQQ13y4NIGlBNf5lX1fTIKXOM4bd7iNFntXm9MrivpKyK/TFwi9m0
qbhFFv89mg2O+gOHnEIHfIrNb+LGvNpeDB/V1Wo9WttCQy3ap1fnao0ArhTjulbGwYV63Ulm2qyY
slrjJiNL/PRPiIBVvF3MCYz6g08+lvDKm5wfvoFY2xn5GxNuSZdtz/83d8XK+t9NjlgU1rNSWdfE
CCD5/YxbA9oU81MjqTDdvmUzf0eX4+p6aKru5vVcc2OgbTT+CAW2YQvqggSTZOu2Str/tLX/gFQ/
1VC37y50lvglF8+TeV4cV1gvQhrdw0wtxckVdEWWyYvsUR0nUC+2M5CzaefmEPJuvNuTlZcHVjvz
V6P9tmShwLEVYS0PbpsfIeACZ+N3j4ER4kpNfhGkTX/pPfLyz+4gzlKEWzspuUeb3vdddXiOa/iW
4x1Q/8QkXHvOEdnbAcE8yyP2U6LSWA5kxV0yWEDIYiqLM0yxUmeDMoXdAHgHqSM+5SP5PldrSc7M
9DI6SpZMVKT505444qn2K36qIjRCGV5kftErrK6OtnMucKlzgiVnCrwmYJ2/cuQMTD9eorU3ITuR
oH3K7/3ze3Nd9R+W2c3WD56sQiC2UmTQMagPidKD3oTjtpegSLvEzm7l9psRGxRuQG8kdQoocwnL
+E5ssBJ28a44J2G0zOCyh5j8D6qiuTVC6IE3Z+5P8fbr2ZvpL5PlrAFRn+zHWztkpvyihYi6H392
AYZsKbBxutsPEZefPIuUZf2heUGVn9Kj9oal2W6yS24yw8YaBZcpPthOJDD8DDlige7bYBnIh3zk
1Fu41FTa891tf+eOTCvOnz4x2Iwnhc7BQk7ySTVkYazA5KhL9SOXOkyonK9Gz3rIVg1PaFdoxs2D
Cdex/aR1i1F48amu6TQiF0fkkdRlf1Bxll4YSPcDbjZLQ8UrUkubVcu+XgrYxqNWAa0G/FeUIXjD
uzgysTLsI7dZwxCh7+jEwT4tkad3ZAOECuhJ6sIMi8vU4vpi74Htdb0akVvWaB1r4f1pyZSF88P1
IJ6GBltMQ25DKb/fVe0pqgzh/bV6kZi8yAGrqf4iRXF1rJ5TsR4KmOTloW7r9JHjAra4mVsTvjRl
Emqr0MyTZQMbThv6yU2QtvBB7qWsxuAoEiyT9EZ4ARU/1r76uXSUHABqPlh307XwA845H2+O74UG
kfAZboio6zMgcPTxm1nYoNGQCzAdZIyMLu9solNeRrKctHnzU+D29iKtt11z3yJ62/3lZbxL0wJG
yVY26pyIIR1pfK0Nti6ww+rm2T2qgh1YMuez8bbGiakXJidILCtQO3x96fzAh7j7Yi7RA6mMRw1c
K9VnDU1szCFgMJr5gI8ILByjmYbeWmUp3Ll0aFB9zvQpZOTxD5OTWoE+YKG1bQO8J7B9hHyqdOoZ
QlDRf+4zq3R6W7xA9xnD11dXdbfTZkthskFfiCi8D5N60hEDiZjbRaderwVzl71F6+vu0S8eddC8
ZmgVPVijMIOYrPHgRMsduzFPXJcuNt3zUzdvYucoNPM49iVtZhoIlnD2ZwH3LJgBJKn3Mjkl8pGM
DAIAnEEcA1hybeZcGySHwJDxV1yg+1y7dP/ujVHy/vWiyH4wC2rV2i+Hg6Ztc/I7lB1D5qwaEwOw
yJUQwsLxvBofcbCC2iNRDhMeqf6/LLqb64v8a2v1qhij/jXFMs9i3DHgtxM4bevIjpALuBkzeFxh
40jhMJJo+TBwjYuP1s/YBkr8QiL5y0rEE+dysnKmt1Pi4j+r7YT1tcYhAydE0jPQo11GLoPM8bOY
cDjFFP0hahuchQcvYOCh3VWDvRv0Zj/brLWn/KjfV/aEhnzs91tUOdVs+KjGaIxj9EAPQll1KfLG
P3AYkWkQMkyLt25osLLtTfB1SZx3LsxNiyxQTCoXBvk89ADLWbD87vV9u0pHkyI28xhvKTleXVcW
88bTwgKQCK98agE0u1+DFeeOWye89Nqfd1J0NDKBOuGdkwqu+jAez4eesHZT8O4X1gxJfqgzwXjY
d4kf+0nvt14Z3gFj8pUZlX0R6htbmzkXCi3/tSNIc4DH3ccYT6er6LL73Kqa4zpRvFcL9bX0xqgd
mOUjrY0M9lXtqvGdt3kRZiE0cu11F7geNKEN20qt5IEw3CQMSqheCQfezA3zU28tRFGuIWO7cYXV
ggUBkYnw/66ZK6yIxIn7htfz8lcAOTep43p7r7fO84oI9BcD+GLoTzsqsYSRcV51xraJLlcPGhAj
JPmkBvGxJ10pqpCa5NJjfOPOJFKiJvWDcw6Bnujv/AI+2veAJfqAdz60EZPqnvRUHdD9veb/o7G6
SrgIZiS/TIVVY4pIX0i/Sp/HyYKRrOMuKSm4XbCiqkkLSH5m6/9eRMhALu2sihZ3QfIfBD6/Ot9u
j9xj5FnuE6/IA5TSaz3HefEsymCLy//ANmlaWp4uG07LgYbBp18Jg44ECkuUd5/MsxhStH1vx92X
szogU46UtoWidpZbZY+XVfMl0S3IaVzwWU/IglQoRKBs0/LpENh/DagYsxG28OvZmIUsCPoc3CVZ
uq28GkvDe9VVysmMVJ5Dn3eZUyqPGSlcHarG0O8nxlAFfnJUJIK80b5q1F2nOdAdCreylzoPLCPK
VyIMeiWUH7JA4n+N6Gp13F+PIjgbKYJjX3vUzz8tdBCcqOV6nhe2A33a5Q5qR64AED0GW5OjTqZy
7tUA0HTuDfM0gX3NO/XMaNStkoNAbyP7mrJo6ogywAAJ1BluMqzClngIqkyioVPaj9kHKMj7LTYM
hwwy4srMjwZkzvjVnzddDUUee5d06crGnwcuZBD9vlrEAJSMRPI9C/KsISi7tO1o/6ei6YdZphsk
I5q0l1hgD4acDoKEhehAsSAG6UVcJ/dDGZp1Qxdw3y9au0QVTPi/JnYFM+zUGdsbO3k7GO3yhZrK
ujAStKfZAYixtFYicMIaU6PfOb58WwBOllSrfM/FhjqEHI3PLVEZ6v31Yhfd2abqKN+tW0Fq6F7I
94HRLXb/Upg9iB5xsryspYHnyjGzipzy60Nz2g45iS9IOpopeSns3Jd+KvVHWeVvHt5SUKSyaNN5
2ziMsC1OhXSqgcQdwXFfKU2Egl7MAf1UOUMc3sGCk6KqmiMuTQPKkVdBmeQMHKeVn8Nle8ojKZhB
IVjg6SguPnJECXMJMo5DTnAmMANWOT8qq8w0ha0kzYcFik8TwMYvOxeZ7gxfGIf9ZmYHVBIhV9Ab
PWN8fdbv4W2GDLMp7JAseeStD8RkxtjDmRwEMgPX8WCaLDWBrAx9oMM12kOFugN5zAoixFhIdpPz
jR73PUr8M8sPQzNQhHyyHIpymgLpiIksgjnKuwAl4jojb8koJeyPcAWNoO8O7yJzYmL+4o8yoU+z
yrkDiPmQ7VIj06IYdr2eOFL3Sb6h1858VjH6nYN2EvYOWaBILTs0Kk/ceJMr5/6NrDZN+1QMlGWW
F8n78g98czD7oZ1jd1xCa8Pat8qu2fMgqF2wuoJhf1ZMihY2hEGARUUW9Kp+tDcXJrBC9w9WDr/6
BnqF9d1LIRpOdGO9viLF1X3W//X2S/gfFPZBZQM94L2DPUg1R1bIcHMd2nZyhndj8l/ZfkO3iWWb
AQctrTDfTn5cMufz6NacdGu3Log3zGfHO2JkWps2n/5O0L/Pgtj8zrCaG8mE3B6S/dynRkmTscxE
Wm9Y1KU42WyiqB+3VQ7Ej4j1KHjYxGqJZukusiexd1tfielcEK36B3LThI0d4a7NTBfEaXxE1XFa
rSgi2BB+V7X5kukDS3w6F2xYK5wtNeO/bAWljT+1Bq7Ot6ormFzWaCdnQOWFAzTTWczLVM2taVb1
bMTg/xo9SQKpTZg8jkcE6QYul7cpVxjOFAYGkTcluYeGFEWoz1Wx6luhThsQAcA3GluKTDLZOHDj
R3zZyNp+J+fU+rMRrche45b5xlbcQyK8Z/ipARZhpaoxw6iSNKynMscJs0hmCmK/4d4g/MD7wa1P
vAFyZhj9FStUpGKvYGHKKHQeZHQVQb/1KDPD9p+9kyCgWssiF8ljECl8i7XlE/hOmMn2rRIcSAAt
4OACobLSCV+YY8KvXbfg8WTwXXHDIk4XCi7SvSK6VX9K3f8+U6bXzOh2siYX3iFxh/Qoear6x+Q1
SXzge65hUs96lCVPF++8+L2c0ZfYoFvxUna2GmH/eJP+B34zyrUd6/D+EYE5rA4mrkMT6vPGlQrk
mGynjGKGp8fV9bYaDXPVbTRImo8hhb5zQlW/ICQNqhN/YVvFjMS/kd99K8lqsJ2D6D2g5PLE1n0U
bbEHtEshv0cXrdw4d53MDXhoLT2lRO4m5MHulmM0cNsrMecIfaMImtCQfN7THPweqZN4M3cjtwuN
Uz/KoHMz2JKbE+BqqNI1rVQt0samost9KMQzN2uNPJM+1Mrf4abjxVyHStX+679tpqAvt7EbWor1
AfSoM3+8KIiH2dPyo9uqDjWEo8qZz6s81y6eekNmovM3D0B6S8Xbv62lggg/VEU7VWwIkXC3minb
Q5SRQudS7JRy5AByUUVycYbOp1yASnD9vTADlVN3FJjNh7NUvkgP3R5oHlNcKBQxLzQm5O6eAE0q
bWSyZo6Bx20j7+HC8IsYwMVq8NIdh/SpGk0fYRJpflTD9KyZf6fteYyJT7FxryRcJvXH++dX7Jbq
vlkTaarqqDoj4K6EovIU9GY9jk6BDV0ZF9pd1fYnpFbl0w9WF0TbXVUrJ606zCPRqpGPWgT+oRmZ
L2AUaCAUXy/sCZYJbjTgtyHAoiTtTX1en9KOehSoSsBg1U6RcxknogSuwFj6RV4ciCgX5EG6WpXP
HUxX86WHII70jk5ARWfIqDa0y80mdXuCs2Q63dyQxDodQ69TiR4V8Lv7fqxvAo34bzHOzuP7TSpt
6kYvIz2ky1lNya9p2P5bg2ud6xzdr3+zQhMAf8Wxl3/RcWRat+7YK03q58Q3DIoSs42mY4FNqkXH
LA2Vi+/L2U+75x5Vi5s2kbJbm6yIB6rLDgawKUyGHJgRU3kH/STb41CvVZz0ASX4mdCbSYGdmZSG
yYO86qdS4bRPcVNNos/o3CyzYDa3KBHYBCkf6/UF62iRh0lhLa67VN+dCZDMDqFueo2kM9n2HfD+
QoczzhJ28669KTq496rY0jngbRd1RQ5zzQiW4SmlMykAhFdikpsZjB7CU9acL6qGN87ZPSNdTW3k
HYdh6wMvWs7bY4PHN52iVcFdKi04zq9dvWUcVLriMeOQNP5s/2GLhoUehOuWrPtLgXb8yG6D8oMH
+rUaWEbBcBbuFROaIqMixZ/4joyNFaFjtK/0CGG1ukLai/T9qHGVsrWo+Qjvn7D5x058C4VB0CQb
Ey6XmBCY16P+4ckMm0sl2QoK8iFs8w03F3dl+OkSvtGykH1aChs75SmGOeX+XbCmIM7Cy3rbt6LY
Kmbt4WorrLfW0mA2W0euscNoDm5FAbk5HRZOA76wv+LT17gC97Ssnekq8Z/pF8hOuTXLCtR0wHx+
iZoaVcJ+acXYvQMKxDJs67v/r9Xmh+BL4jViTznugz8jC/9HDTpBqsYHHgPyJcbMD9oMcIAhAxuA
Vy74q6rIxV9BU6CXB/IKK9FF61FPVvD+mT0CMxRffRTwQERlWApL/SgC6tc/Zy7oINk0pk5a1UA+
IUAt1B1/2Tnn4XGkCR7LZHBd0itCXApQPa70j4c2oMJ1EOot/+0ATTBJh9p1qf47Wl3APTVALbsr
6oJ37N4zak8OJgnqkNaT8kuA5kUTQSDvxacoNio9c6mRfx20lKmSW+CJqv3xOYKL3XkM20CKXtSD
i2wD4ZnpcFue5oO8H15d8V+7EbdFWXNSb9AS2qIZ8Ow6F6vrAWH5W2RcycUHhOBdq7JhHWZjpkdV
G9/eW6jJQop9opOWcOCNsm3oT6wxbQcvo/bPRZJokMSKY7xYH+cBecZfSQm+47n0RVv6mVtAuPKS
SgPCc7yNKPOBziGHQiLh5fFOef7IdjcMfpvc6uPSJpD+8ZP4f9E6fzVYDfbzuKCp9GW6uvCmky8U
DC4UQ1h+4fa25SpY8fsNzp9xHAN93DlEpxZIqmHEgUsYYR+rRGF4a5jBmJixu7Oh90KlRLk9mVbv
ybDMHoj9zyxYe2INFUxK2ljySGMbp/ejcesHQhrgdW9/8/KwU+mOpL5sSjF055LkNC43sd3fx+r6
zpojb6uCYIGjxJ6E1rDzIB056h3ikVvkOLKy6h8AI9xIypDODm4jzcuRzFhp7YXlHgj3ymhgXQjh
mhhf19FJWV4SHPJdytuv1GARDnci20/b/5b+2EGNYfRb/xk2YmO9GjRltdVStFet1CoI2arYV8a/
mNHVhdEfGCGtrfKakt/ckpT1OtnYHY40wpGALCVcRn+eQsIRIj3qSI2RAyiG8n1SaMcwRLI8l2Hc
R8D/3k+J7GN0OygGrcohj22pQIEnlhWCVjljyJE/5/ArQ+s+IyZ4mumM9FGdc0whhPfALq+eyq7w
f+kzUahQ+rx233sBAIkQq0K1pogkDm0tSVUJaEoA3+uN3q0cqijpTL+mpIH+l6578Y2HhCgLJDKS
/RGVEs96uG0bkK0ymmwFDa4Q8Fi/eLcMogBqDGEkeeublNo9JkyNrYMqil7yNfeZ07QpnQZwyGq0
WzvHzWgfLS0kOBOmkyyKfVXduThi7ek2eGDKIItCktZW05KNEBK4ZJW1+Lw5WsTLgBdKZ/rXk4zG
6/SUgI50f9KNxvqC8Dryb+IAKbCrurhiU9j5P/de36izewPcSWVYtsYKby3asOXh02zyZXJuJTjS
9c7FBkbKkCTmMyjmpODh1vYmFyRdJNGlVkrzi1vf9SBvaedqm7WgXenFnsdJNgPH60IU1vXWujiS
r1qcScZdcHqcjNlGNnioslpswKH38ZAgkpsVxP51lZk89CkxyuCWLYLHj0WQUkJXZ6qaqPVhOfu+
G0Dql6+Uh95cS0lwjRmUMZlV1JIsrhEWdXsTd14kWH7/BwP+QOK8HSGw/Ez+sKjU3HbtqdQW7hGX
Rzvc/Gk6LNjRW4vTxcN8NwPTXQbFdhnUlGSAbO6lrgjgBUmND/0INfCqIiTCX9PN6lGoYEvoEfE2
eZ96bFDldMjcMA540Cf5BpsLMmUkF0jyc+sQgpJWLOQdiveZxyn9zuejIGQBI/ek5XpYn6Ry4Xcz
8C3ZaIm5SWpV/3xyxF5XumfSxVihrrFzp2tVN+Z5BcUxV6cGuKANgG/Km5EHtuyshGBnCipz4n9k
fsn4UZSx1+6+bTONwXPqy/RNCAG5710RtOLTfhiQjuNbJeGvEBhW85R5tGxbakwM3n7y61Kxob72
eEHU+WllO1XEah/iBbau1xqSKwflpTuX+qEZzgO5p2grHvynyekfhpHvHoLT2YepDTJHy//yUUdN
JP8ynuap4YC2C9gJXb4q+jfungYe2XqA8CuFgeq9oksZ+WCawk5ktBZRz0OH9xscyVa6XAmTxNLM
grz4R1GQXBy5EIIwmooBO9/pFlOMfJoPz1wPQQZlfqOawgoKUOYLrnlyy2wp3mQHMU0qL/bxyLzk
R88SaXXAhwv5HAxmnwY5MT0Si9i+S/sv3o+xsoyQlt2F0qty+IY3ySiJRUN+6JDtkjnAkuUxnlNl
hcQMxX3GfL0CXhlHjOOLe2h5JG0vFWyuBKB6cyHVG/x9e+6sIDlUrfkI+ZUxm7804iHEwvhFYeVP
v8YiNFTwNWYh5JFtzD72zRol273Xow4naFm9KNiahHSWSq37xPWFUmm4f8inDmoPI93I8b0ibKsT
Ve4Ow/WFH13TLDINGnpdRLZkQJNScwZg0yyL3x7cs4xhb6deP9PtTyMo4xVqq7Ho+zjPVkXZGnOy
dWJvf8wzS5czt+45R0i2lYymKUkr78XsR5rWxxQcw9cDCEETILokT/8QNHgD6jOOXRU1D5dX2C00
cqfnlIvCGf262rm8h38qJDmqMrJbPgvcXxY7JGxrv6mGN62EtjNqo2+jSH3IH57yRD/bo5yRBCAf
O7g3kmjvwLNYUtl9g6tbrsZ0VMDf7XzGks5NH7OYxqUfbgks4hdKCVLS8FL/7sqH33zc/nsFMZiO
0bzLwZ54ALUeQcP9re6eI2PnOiPB+WAPiURSKHYVRZrcwqiXmse6zmtu0xSNQRadYpE5WtE2Cq/K
XtZjsORNcRvgoovyA5cjQC7JZer+e2N+8lkbNQ+r3rpRkfeE+qoi5lW3nebddD4pty4o32MJ7BoD
uVlJBBztIDvBEzV+hhO6RjDqw5aNOiBAws1FcQQdeW7WocGuIbRoLZnOk/SjoHtfBaaFh0DsNmfJ
pegjx0wriQ3knk7gCNdJp7tSdbGWRT987XC8JxsVsKNKRs2z1okMbzjCc3FiQMh1n9L14wQYb4ei
eVOVhXhd/qu3uWIhWIoiiHTVNIrVKTCk3IxbbWM7W02uhN+HYFtJs31bWCo0ipTiD3iSm8GU1c0O
CnX4IBCZrursZVQWMhfR9dqp8CUfKwTkLbZ8/pMzFZuVmYe26c1FS+0H+fOWPkzcC69EG0yCR/Gi
+mYty+7oKVZEr0c4JicgOT6qUpBTBnBkCn9pOd79adtilnd0+D/ACk+EOV7qKlTulHWMyM8hfl3t
l/wQrKTFNqqbgLWcycZkPk7Nha2sOVs9VZ1CIJsmCEWKa5LgoMMQ+o1VCh3jrOklo1u8vUKpsrXC
AoMym/MPH0JhYdHF7c/S6/Fg0w59KNUIGUQ3ufIme+OpIpRhb1oBUYp1uczlYUd37jRJ4h8WpAVo
Ai/IuykYaZ7aYZreunVUjea803Ggnah5CzSUoUoIL0cSlH9xyGbnwBJRJFs2Bae8PiG+cyFMJda9
eC2fw4YK9qGh/1hVBBnCHAGxKIVBySKFNLWUGLwibuCsYl/xFLwiICfThZWaDQHa0P0sImrvotuL
yc0h4CnvlGdZSjKNiOomJy5A0F0MTa17pDuhuwTVNhWQDL7HNp9642L7VubwvWU9gLg8w2sbztvL
QZ60kIuo+OzXb9QdKrbcSq+5EFreU5mQ0KpkfCAbm8CiXvX07WLRftgA+KqFjxaRhvi79U2yuswK
BjTVszWeAQ+ct7LGxwJjztUMCM/Zdq0+Ei6yKC1U7raXdK4PL7kFGZdHQWplIO3U1h/T1j+a0bgY
lL4Tan7iVaNhZoLQu5bN4KfFPgxlZraIgxjwcmx2l0ntuKAYmG1qyTixIbSxv6ZnBvu+nOomPGGT
aAoGVkuLLbvpG+nQFeU6lz1RLlwwo21TiJl345ObVeVeaX1ffJzioDP9SzXOiwWmT7RYHXTmFk4R
wPVFV+OeJbD2Yj+hLf/msuPXBXj6/YsHWxEbHz6CIiUA0WJDVVsKm1G6J5cFk4aNGRDl3MmNGFF0
LBKAZZTH9zG+JMSC1672AjHAvH1NmAj5oqA8VUgKx4KslD36fDUEErVzQpLzygfRfs4Vp0pcmhlO
LITOwJDvDseXOOwoF+ubORKqtOgSdrNDzUq+kf2nJ3PjYwX9QAKYxHY0o0qBgdDGw0G56YV7CBi+
G2QeVSZahsmlr+0Q0kwyzS2W3AiaocH5adxrMlfWnIe5uuqTzy0xo4CMjcITuR1t4cm+ApzU8CQd
J92fF0DrVPmf6O5WcKNQYTF16Ov3y/ZRtkF0qBfeinpKDjsGbzhyKIYJXbLuZTAwg4Ts/mOE3AhL
AQ0zjsA3EUZO9OHgLGtCw0qRDVB3cSGJN9rCddgST2MJ3Dijnglly1jXdbtBP+DdNIt0g8Ck4sy6
/R6al1uSVJ3GUC4f22jqXzQwR/+8P48VB6SwT04DcQKjCH/ly7MHKfVsZPAqGL3gQ+gqFJHcdiIB
4UI5+dVXsOxVXHIPkqV/ONlfEge7jtrJfYteRyY1qVzWGrV0WcrySdDCV6BKGGc/e8g1A1QmvGA7
7lAvEdZAYigTA8x1ag/BtYsobapED7pTcVBXAjkqpe5YvHPWzCwcvHKjX7tvuEZAFyaoACBL6mVc
cImXyLHhgg3v37prvcEVjQnuhp8smfS5+D4NcwE2VwrvbCEe39aK1q0DX3sGWAdhvlk4sedD+79q
8ilTbhHSykIVtrVT5eyxS0aYpH6qderFwBUcTZJ8CY9LgWiZO1EwUkgirKBaFTYpce2LzqYKO58z
BJWGdboOKvvt0HX09zToQqPqqaVAMFPaTzs3RELxnhihixjEeYlFDyehdJPCkFkblbvKt9Q3YNdP
nttVXP8zgMi+SGnuluBHkKDTvuUFCegaBFMz0yH4cG5AAtaJyia+6gm68iZFnldDw6yKIlED7A6H
TD8ucsKCY17bcwtpSXlTyK4Aj0JCQHvYeq2is47w5BYo+fd9NyVgaZJ9vDXSfQUvvlZp7dKHoOd6
/oTtVMdX70gRm2+x6l71PR3QJdNlcwyS0WLLVryYLnuIFA2iVvzbyDlVym9at80Wnw4EapibnExt
HI4A0EUuSIWMeZfiv1METZV/z56/S9oF4Rh4uHP+vFIUajJmy8WMHUfX7Pyjhod4PbUTzRUsZdTV
7GULNybqeifXouATi3FdKeF8wsqO4zt6LgxvoCt9DpvusgzcssPLYxbyG1VHog2ArR17+AhTdcPE
LD6PKJwnvmpKugk8AKsvdut1oe07Y6QIjy5pSUye38l0K67jbbNv/vzxw69Azec2hmAcdWgnBg5g
dSJPMV3sHbPexlrfVBCdcp98Lt00kUwSeOV10VIGaJr8suiXYnOCJO/eBhKIsIblki8KLXnmkfen
O+n6l3M+bHNa7+pSbapx2eUYQNuuiOITgO6BMUBB+Vp3Ww27FqJZW2vEttZE0hcV6DiX/6NZeWfU
dQLkNUAw82RZEa/eK+MGrvZZ0XU0glFdMwvdymFgPGn1VxXKchVBGFplIqzSwzIMD6slkO6mdJy3
vsksfaVCsx4on4Ia4NEeg9T9Q51eYiTTBOpNlNZARfD5kJD6rC7OV6J5kpMxSxSgzoNbKw99XZBX
DFIeDx3jM24OrQszhSxcTdyh2WnUlaUxC2lKdFQiQIUyLKT4vGZqKJTLRv0ctbcaGTr8/ZKL7X9X
vESRRSVlCiZmGln777zjMCNxSSjUqDqpNqNs38RDD73nYt6l68N0XNY5U+rug1x5kSTfkT4jQpiS
Lt0zQLN6gBphBo23OzrASy0fm6dT2J5DgXJ4MRdw7HrH2ptxADx0PXSEV4vBOfQv7h6Tu3ggFZtq
O8epENZLce+awjkY5SSij60m9V5ve7h9JQf0M7CgiBI6LwvRIseSOHxF3VkhfynE4CZiLreO4BYR
ofXC/OGwSJ6NIdmCaRxjcoUV6Do6war6LStwinSaWv2tvesSDYHLaNJWCR1YZP0ZFv2IEyvfVzLh
1BxbBGL3RTjHuOBvd8sth8Oh6p79RAmzVvyRa/imNYgazZDw2dA9rqooS4n7w0QAziWZGb3Qqlb5
55kIj2SxymDeMQLpCtiBUzWckdW/jsuzF7kwH2snQ+IGvTyUjYFx4pAhsoLOayPdqNuYqzdqA2pR
p9+XGeJRpC9gsuwp7C53JZBJS+uoP7epSOYgLToE1VEMVHuqjMLh0ZCkGgvdhvHcM3tD9wja3edO
7IyA5XROOpv4ThL5UbZXwIzE1fxC2oQSllYGFYPKrdnxNNA5RGyzLLP0jjszOO/XPGcqFU9GpEuP
B5HEwFpqptOqBdGWOAwBton/bvqKqpPfX16Zjv1I3UD5Qq7uo2QWbRDBWhKtlDqrwq8NzUSU7VGV
L4iJnc1GLZmD/541jLVrWYEieMo+9AeA+ZpsjGBzl9Y4qeLbfXCVQYDvHkJIPjlhkWti9C+eX8Sc
SvI2P6WiCckI27H/SI+SqVIwH7RcCokWrOQvKKpgQFeDRMeb/uMOzlmQMNQr1tHVz9x/rgLdKKN5
JUXcFuiTQV7zOTtU0WiDqBozDCZFpmpueTjeHKVKAjwQDErRBq6S0KxWfihGoYQ2iUce2//Ca4hq
/jr2fMnHe3MWVzqGhOAizGxPWiQVD9yYwdeKlQm1GX38ChEgKGYLgrCtpQ28D7BQj6jk0pOVJb/a
tCUL1HVsbg/awuEpBFQyZRvsrjIAFSAENJPZInpJKOj+gQJ031KzZVxzVtVK6qAn2+rMc0hwdrx4
G9rXOJdP8Q3rehproCKHJMqls9aeaDqIUZGczDps97GhRfaLcTMha3eUxKucHfagfy07uL2kaNwJ
fvaywdk30p9yKtxsGc/znv1fQDrm5L9Bmf/8UVF4VnmUGRDNRixgD7m9yLuL9cZaUDZpiOdZWn3d
Cs6S/fZeOiRYNPzugMroHHP4gVKsa3n4wWEAZKXX3yHnWB/5vCVtAZt5/9XvI0n8CEnqnEyzL0Vf
esGRahLNDONwhDi2Rrs05uH/AzfzOrT/qRtnj0rWoxMMuJm2++cKcEjXn1wf4rykwpn6JvxngHa2
gJ+x3bfHSGBZ1uxF3HKG+08+Q9lAHYUepRX+dTXNN0mbHk8ozNkKsfk9s40kPdKLUUeceRqe8oov
DUB5fq7SosvJXpFH1MjUCgNsDH7h7lMim8cp3zEFnBfAJ7DUrmd53n+1/y+DELd80rKhBo9DOwgo
jJwgeHaMsDvqkq0uDhdd9C7a4NYVIgLPHY8IaqAxsJQzbfk00kFhNutp8WybQzwSBW42CgTSdIfL
2D7UtOJF7Hh9x/w8q+8C26cN10mW7Hbazuaxa9X21dL4yR1caoe4HbRtnJfOqgcAXThTmUrsl2l3
ivLkUitsZ3eANdf4vuPSMXBcx076UHwKS/6b9RR8RXGxJyH0HodoR0G+G0AbDSs9JJr+BbthgmG0
bTo2qV1JRbxKknqfq2XsoewPAf11lmraL4/Rj4nEnAtE6nE5yD6Gt56TJ9E2XX3y3NogR5xNWCoo
7fDEcyGvh3FZN1GOp2C89/JQaPF3ZlvGGzI8wHz1Pq0qB6iUZ2vRhZxlpucvk8FYZBhgWWSAves1
u6bMUKEvxhXQZUenxkDoLbOYUr58Mxs8SZkqKGE5WP0YqmBOMCeYQsaeuU3LgoFhJER+YfM8nvdI
dpOTS1U6Ii65Lq5HMmi5j64kyejm5Og2lzvUJ/YVBm1RpzvSUuwz5tge3o1LhcSAJgqkG7sNsR4w
JHuAAtpGpRljhIQfYP9tb+ZMJhTum/MN2Yatd/8NR1J8nZD9+Clkuuqdh5gEuUhVfdPl3VNbYq6j
D2lv0bTYk0qH+YRz/P6go0BoI7eIjOPlBkN667k/1AM707Z5SE9SSivV64+0a/PmCl8ur+g2Yf52
DGcROAae3Ro+mqJUcCAY47G8mQLIRHJBQwTf4XxwyzMBY7OeBX5j7XTFKaDVf8DvAHeanBGdpL05
XaWxB2Gc4FzJLAoFG72RFM1ACvKcA82zQKvGKVQ9xL9Ka+HI9yLterCjB1slENCXUJTkVgT5emWk
b1Vri+kZ+HXgH1g5+5wLqfmgQz9KVvbUTPOIZOu23Xpm3me2sHraZbzuA46GXOmUyT5VUcQMJPCo
gWl0fmgtmp2eTHVjkLTSRM4uk+wSkHxmtvVvc3lAnsUsYMKQRILeB84QgvveAZmBFFm2fREQLS1U
l1v7a2FjwXiKIV1TNMftDr/X+t4XwF+vAGCaTsDpRD4Poe478fJOK6EsG31XO93LDBCV9gsjDK9h
eGUKr/kUG+P5hKUOueLuUemKg6qOMiMjOUJNDF5mYB1gDSndFm1SsSo1rtC0tIaq2eTr87J9gIlT
+1bghtrYCJJ3aKa2fzAFyhJaGwbjTQd9vey0GFveNSpTda5sBFfTpdCpFO0zIEcT2xKMnU4kt3Dr
iMn/p76/QIT5wKVvEknDzh93iwbkeddBSoOPp6+s/YaUYqjbpTwOxVKvCUlAkumhJWXukUQ+4XuE
DBji1V+KmGhLKHL+nDL9LqK0mDEhKfFgEvVTxyevPANlGRct75nmVQ+lbysTYPwNecT6oSWBf7Rb
BmEvpGypRyDoykq0Ds6r1QYi2JaYkmFOF2nEoT/4w6z5qPK3pcVqqjfTDwl+C64FyVRrt4nu2Aho
wjdoDjk7ol79iTcfih000yH907CnagDXDazkTxerV7XG39qKCaMPahKnnFA0KN23ERLQm4ar0ktF
BrHzBk6WEe4zxGew4dfR5rlHcAAFU8UBTpQCl6n6kpuvfaZI7SSB875jw79HmowYRzK4xD5AC6RV
FjKoPinF1X4DTkFPtYCJ3zh6l82L8QQqduACF/OhZcxpL6zkhrqsC0Jpo/Hnt+hiOAdTwsulJ3/d
ljGVX+v7JlNa9a2mlZEHRsPDgOJvMHKDPBrLSvIsMtFcm98p31lOsyhstDUiJ6I53UQ7kYOBgvnN
S7TALn82v0svY2CCCvwU9ubsVIYj088GUheg/Emlg1+TfwuZxioJBJt5Y+s6GPUwD0lDjyu+eKBK
1yMAIb0zQenDRbopGOE7dduMvQnseAAOQVWysWg0Eynszzq2Huxi899lIQmHMXfS8icdBuYYtGVa
b/h4EL1Y/k4wNRoni3yOkHXo1LSWqmmLz53xQNLyJAjHM8Dkgc7upNVYeVKt8sKOKsexar8CFeCb
mbRuXzEq48zxGzBGlajWpNheq+3YyoYFVK1Ya8DS4n2sMq8TXEJlHzIC7Qfd1E1DonDHmDN4GLgL
gx18kDGHcuj/DPaLZNLZisJsZWj1xKeQZaozLAZi+CdBK7vbPXiifb+nlqC+8pT1G+944ydBUrLH
Af81oiCyoPo/Wuy5jArTsz4ESiDWW9EmOTc0x/2WmR5+5Pv+uYLDTthB5wHsFog8Evt9hQkg02Wb
ahgvvNI0UmP+zIumG6l/cEtwA4PUaLKS5L7egx01cA71V94JmIj78Eci3H2NDYdyzFt1Pa2UKPrb
wYckblb11CfE81Z33X5BraHGniCW+WI5v+zeSaDGNzqN1O66r+R64Z/J7QE4IvZtiVhLn14+bd7O
NDCJizh61kJR4FOZM871ebyzVwUksNx9ZWBUcMm5qNpoSk+afIEZ3p5rzTxv6+Tp5gkcXVzlaTvv
0cenKzkcbyYaZ8tmsK3eR/Jvqy6/gzgCn7vGHxPega7JW6tZjuF2/SYzwtIxbpjmyCrQ5Sb3xykP
Ijk56oMV0gaCQ4RQyQYvshLvMuR99MA/AKPhMTEZeEWvCOO6NQ9cwUMwklK4WYXHKaaiAuA4iMEf
yAvec2m+MsD3p9FVj4Z7rsC0++ULIlRz3Y1QUVJ7osYge74bzWdVYog4IIyD1gpnB3IJ6mcdkplu
jbmtID3GY4HrXgpCGimEXBfQOCSTKTWteAImsIdplNq5KW2iO6j0Fh5b/+6vLHD4nv0k+ArHWzz1
4VCh0mG66aDJLaNQhJVj805+rChp+QurZVOLOFW/H0z1kodN80Qu4kcaYm5lmZBLp2T7IRl2FpSz
K6LSOa/Slm31oHXFJHi8L9n0lCCN5J9KBhts7tRm1l+5sA8k+6cit1TXcm3rzAG6RB4hUXm5ewar
xpN+1f5EnB6yGfRZS7WlUP9svHqoG7intzBUlBJEYLQSlKfRxzhe29JbO/tv1dg4ZKXscbiXV6fh
QHNOaP4cC0VELBx+nZY2jEb/00SCg7GsAMt/N0PyH+ohhmeqj/fUksgJaphGd9I1o7R2RFMiRtDG
oltUGNkVMoYNvP9dQTJstJ0FygPtLiM48jJXNR2+QltJN+vsPmNL7WLKCiJP62lKtd1QPw3msWA0
AeFTJsrCfl8jvd+spYljAmzkDf565xXWh4sw50VgVRa2MEU/knG+IkqLHsCBlsOvoqVf9HltU0oy
JcKfvvGP/gQcYqHQfitsiIy0h2o70X7BN3jkUtdAjcDDudMHsVYEp52uDPP7UgatoPALQtLl9WEu
nxN9wCnCUhDYoV/Jf8rj3M7IHepdSlcdt7MrRa9Fmx2GgEiPTFsWONJUge4redqH0bFZZEc+mNBD
RQ0KbVO/9xK5qgkwzIqrpa5pbDkIqTgjONfCKvJEjrybW1VZ7TTKhNeDfDAxnr8UvIWqaYSJNaYW
bEeZER3etc3SofaUiSp3oml0OMEr81xYXbTw+Huhz55i3+JV3HbS/6zNn8LMMT8TdAmA7egwE7Ny
vW2zc1Js4bM/fMab9uHGqegGa4fpj1y7NOHg0j5KB4yPjfObeBAXe3P4Z7DrUMk6Zt2uLlNgTt39
/okTszWlkU7UTFYqfVR72dmEEvt3x+bybHS8jnePoX0nWXFqlr99mXsWJ4BJfmU4Sq6xy2ECc+4z
rV8s6lQmHC1Lz1904JXWRnUQFK8ho3fZUq2jKzKZKV6/V+Po4U1Iy6svAgr+g2vcKPD//SsyCzgS
Hvbs1o59wfbOxu7I5G9mVAhgMrut/7QG2nBuoBWWx9GJS6AE9sD/pW/G/NZd9zi8pbw6pkYwQUUZ
SQQoTfD6rkZfSFpJvFXKqAHshjBf9Lv7I4T9J+V109eC9Ed+b6LKmBb/roLYlCzPEI+F/KW46G81
WXrch78j9quH2kqqiGfT7aV9cLXNUi6BQwOlPXvCxjXnjzA2N4jc5aRebDt/q00hKHhhFLpFE0n1
JY1gboxQoshZMBCrl17wb1vnxrYNUt02ID1S3RGkZXVLeo/r/rH03PMpGYiBOMjXjhXZjYXsJuwM
a8VaMeU5hOwBDHNTeB3rEiuYU1b/XTozOKhaTNtlr4PlfeDtplXdL4BV97Hh8Zz/Z1gff1YoqBdJ
E30TvX3ql0CCK5+WpEtP9aJCo417PwbLypUXt7DTHMftiQp/DUlIGU8rJgnWxJ/mD9DFR5Tuj69a
bqV5Ge9Hi0rFdJbsaajbjoT5qxc5fIgnJBKzhfI6JXU/xI1Wdz8kXiVLMR1uL3pZvxoci93Q78b5
OGCC56WMrXQCDc0TTrTlztMwsTweMAbG1dVLA8lFRh2dQf92AsutJR1K2QwsQUo3KKs69fR81x4a
uqkG0r2h/l+eSkTap3C9rdRKUgK/8A54MssXX9ifDjxkChKcU96KNhgB1j+JlLOLEpdwagdY8uWT
BS2fKAiJzGPn4aY1EHQEEnvppFpmJC+NpNlMfAMIbBujOqz02H0vczVBipUHXl1IkVnSUWc4WUjF
HbZZ5xUN5dQXnPssGluoPULwigQwSl+FA4wIaASnyCZDI7OQqhfMZ4KZyARVcEl3r9Un+4zUwGwL
D9dzbt6d7BWV5YnFPhcF/BRs/RR5jvDdtmlvnZmgvgTrTwCUKykdMit4aDwc/pzS4ZA+tpmwvBtx
F1nXHbMf8ffUlrGDXcJVgvt6vS2RgfWzsRUlDJm2eWMzqCbGsiCzD+KxyBb08XditzbcPKSGt3Wh
uhbdKW6vaKwGoyKms5tj8l3FqY5RBDnF1+/rgJqRwCXqQIi+rtBZXLbLIK7K6wI5eixM2hdAcOmH
rT22ptJUrlnCt8dZxQYj06P+962Tx1G9hTrE/ubxbxiRsBcIg6GVY28Lm1kvW4M3X/42YGN7Y8MZ
C/c2VyARK3TXvcAeL7TLeFNnk+Th7EaBKhCAcuwHq1nM4MpJc4kGStqgjtreFaNDKn4Dd7kdhZcY
YJoLpHcinhLL5yyTzRCg3kdsLabESukWUQwSomhz3xvQZ4h2iYF+LNX7Zwy60y86qscqWnWupGgp
NADKW+QPltyNBOHk0jWvK3LzYpmde9hm/rHPXcTAqdhWfBdC11OMQFR+sP41NMtpwMf89fPeKCnE
GlEAK01cwmQsXQlJb5A57YdzKDKNKMWE4QVotMo+gSZVVTEcN0/hmwOBTp3l+YpVYj+RXQ7A6aYY
Z0GG09LooDd0emXelYoJ8lwupOqjZ8mPNzB/4vw9V+9tb9/eE+Q0Iodtc10Z6GPFufBZZC+vqJIw
tjCSvx6OGslExYX5dcnAlkoeLODl0Vx1fril+1yL7r1j41CVJoBHQOw4o1RwyEewHAa9daRmmZam
1yissOzKj6Aw9rzRrLjOqiU5cjlQ7Jk1QOPw4oYH2MTh1TDzyFIBMhth+ERRWbnk32LQRrE9Jdm9
+++htSZ9gYeDLcniGm7sNz2HspIwF34Qc+kgGRkphYF4GhLyfZJ8WJh3KLbzsb21zRdnaTS5w5ir
LOQXCY5EMTfGul1UPiew+5/swb8K4Le477F43YeCK/qVYlzQSf+3UFC7UKJHN8lSYCDprcEYlr5T
peFUv7qCGVPjf1QiomPWLaXJ+5iq+g29D4DTsB/YOGcfVpEihUUxY6Pjxkdq0eQP96216hYrewMb
7attxyEbYqxMuJ/LqYpFbtZEndP2U69Xlq2DqsOzaCAWhsjxa8MPIg03Tr5HulMJf2zOfAJqLHkA
TDYfBDQHI5zf7GWe6nNx+ptn2oqfbW17yZmFwNwGDDYqTI6B/21UhfhHKQEwmIAU7phi2P+1VCJQ
55zp2DiVL/Er30b04kTSvrxyQtuukTmFggZ4lmyU2gyXa1ek4jx4zDTvQckSKxDCgW/I3Din9ru8
kZ2wKxksTDgUgEhSks2s3IA6UlDIiORViAdj8UfgkBLeM9c3ZSTQ9vNPldSyyK+ik503zDUwXhxn
Oq0SRJbv7ys9rybPC41HzGMSvR48bc8QYxHG4iyP7nwBJiVgrAAnWtaJ1bM7Qi8chnryGoHFZOWu
IIJAfWK2vXvQFnKRwxTCSWYuAA93oeTTExkgiG/7lqb1ClQ0nkpHBdRM4Ws5QHfiDJoZx8tsRxC8
lH0Xm0LQcD231cS2kAZPMk5wqJwl2kK3mJK/p0ODVlgZmVTkUTl26HXSwgiS8P0GakpRdqXCHWnu
+fw5bgiD9qfaC83DmHmELBqErEM1v6IBj3Jt+ad+vpcYB5PM81chMIQ+f+vtA9ciLu5L8fpiuPgA
aAX72zHBI/UMEJv9mlIP99V+1u6M1fk48y1jCOcXbtlhuUjMGfLRAKA4rHafqlRCT2xkBQJs2iL5
yiOK2IV6WOq+uMLiRL/UAe7qh7adrterTTTDk80asuVr7kXjM7ouKgix82+rtbcOnsfihpSZ4nUD
wR/nHnai2vyQqlgwkHFjK4uURK9lRaJwpN2VuP1a6zf5hSBF7CS0mQCcWluRhUeT96NoTP6l7FTw
m8BTh8aF53D5Hw/8oJVKGcfNlVbL41Sod40JAo6UJqf0haKQPXRlTwNZFWr40qKmT/zY3JBKY5k2
N135cJRvtDrewUiysehrIXeBNlKhoze0nlF9ZPfeH45rNIs1KTOMFwkHscDOG/ArPyQ238CbTagH
s0qmtlkCt2hyFBhhLeVrgsufiT70OXorywImsCM6rCOtLpF4NRrQTCz05YRkSdWx9elTdXnS6I+U
NoBN2UfOt+F71rTEem3sjpyhnUz5cDuSu/WNe4zhNN+AmxQooXoq8EOY78b/BOkPoGtrixgN7MDM
IeoVrjeMTM3Gt5FTRRyizZuf6l8n2fpF33d7JR/0L8ka85dX9qaOhr97hHZraoAt0fVrGzERSS5E
vXzxrd45ZTM70GXWjkFzKKNXJckW0fHSksPapgwy1JURpKZZpfGXwtBAXoFHFa7ZeYxJUF41cMdt
zNaVI7TbSg9RxrCNAFyFmLVjdTebysGMpGhsXM9urpd898azcrr0eyG0JiPFP0SL5uKnwcyeCJhu
ZA+NSsCvNzcgJ51TQon2XUUJKK9L/4rkqDGoh3SnNNuHV+/9kzFhGoh3e5ewrlqKO8/4JdaJqhfs
IwpCKPy+DWUCwbVN9kE+2ooaUqjeRuUfPnPZy6bumtC0X1oX5G/uLwbh6seQlUzc+vgecLMM8Ks4
kOJminX2djzWxp/vBTlK0RlTJOssDQyX8s72Gw0OGZC+Od686u66QrgZRdPE1tv5ASukQxDU/4zV
cz1B3OveqWP3pivqFdlXBZDO9hnOGM9/7jn0R35dloPyagtyrGNFg6B85EAXqf9vpZLU/ovaM8ZM
HZiza3k/vwGrwzhr+NJjg/qE2Xp8Q+mKZn/qR+ciqYhs4NIW8ePXL5JFg4Zi+gJldTneI9RIyxgO
BCPIVqZUtqeolRxFlLTMoG766fIArHdchbPr6nNEN7GmP4GGxH91kSCfEvArPB4Uwmybd6upLCbu
30xmzw/sfBjZ7F04TsiLFbGgQ98ZffTBW3uH99HuQKzEiKR5VqBC//a2H1yvI1piDzZfgiYzJxyz
QKhUHguU2EcampRJ0BH0kJSVBlEyp6XdX5tS01rtC+EnRv2vrMechjuxpxY5nqiBKF3cMEQlESCG
DsC1TsNWGQECCDGdsev7zsaaReWOl4pKk0ryYkI6IcsJiLrIsHBu5E+VewXVr5SvJoR6z6Rj0m64
jaKQkAtJfVC0i21sw2ojE4xvwUkyNn4r05IiTEWkEdJ+1GbEluJt9BU3X46IcsaysvxexXBOiUuP
t4HKbum/ytjq2MRLR1hB80jH89Nwra+3vRg5o9YQ40/NGQVkJ1N4wrcxYZXC/ApkAFTc8BFEj8Rn
YuS+QkXcTxKeldysq3CGOR29kDpV2Xchbe6TpsldR+vRlYjbwVVF2a5BFWG5vEpm7UZueGXKzKxA
KCLA4ybYhJ0GXwgSRNP7kNy6Hr/MTb8gPYsblMLcqBX7M43n7jhRDg4qvAI7FZ4KGofw0Vo3trej
NeLM8xPOQQ2Qfenv00eLqRmSo4JFW2mVBOGcfKE7te0ZiI79X+NIdxE/EfnP+3ItQk3dvsmIRi0m
uoGxGBTH4+H+HfO/VvE0P5k0fn7gwFCC4SCWIEAp++Q2akdKIiE22+F6u4CSd75XVYpJjFIpRD9g
wACe+kp+VCYw9CTvm7g5Tru4evlWFRXHdNScHYy0CjFFIjhFxh4ElqD6JLlTBtVmZsuHw3IpnNIj
4MrU12EL855Tj2hokeEfkN+1RnFqxXyd0aHmzxHRKjsb6YT/o2Hq34eH/aPF6gu3j5x86UnfIUtO
9QntDd1FQUy2675A2MEYVNH04fusDjEBPNFQEbP+UsdGNMUAXoFKD5kqClwd/0/up+QTWiwe7TYF
WIcbdJehRq/9PWn0BVzo8jcLB6P1b4j2ENx6keu3CBiXswWxoy6J6+fLTpHpfJJSctA6XuOX2v39
SmoVSfN1G4SPCUGRNO9uPju8YKcylQu3TsuVICRwRFR5oBOWQ1ui6q+etL1M4tnAuB3m1Qz6BB6a
5/cS3yq6O/7wFC/55n2DkbBZHnYq29xDdRWrF/w1hDiTdyXXVfIL/bFYo8HWlx0BsV5IQJzdAvLX
i1VJKDJ6OP3+yWQUrggt2QlFSITSlEuJuLdjm4BpHnzz1VRwfcWVjOB3DB39vMm/txGYoFKzHwht
I6oxPJDKKh49snia+rrUhBIIFKLD/HjJgdM+61WFAzXtzafhvO88zn/wHY6lnRQZUjWJdRgFo13k
rgU+pG6GxMbkdfu/OmOyfsQOzSqJ2A+EV8ZdDSazMB3OES0peHTASU/DdPEKbppYBmoVNCeqLNTP
H1ZF+q4AtMl7r8qmx2/7gQ/BUHQOkhM0ZNYhFT25GIoqZZ09okQhoZJOFAUlBcX3qkmz76VNwMvE
/MlhOWCwRTZdU7dfoYjX+cbS7U803kA78X6aMiL2RxLVY6BZWc2LH7z9H00spyYaCQ0UuWBRQuUR
CQHvqA56v5Cspih7tkJOfZk3WeNfM7zvoEJz/aZOmjEQ+bHYgAYPCpQ4m7KqRdivFEOTXlovXeCs
mvvImu4lzhc+mYtX/QlhqA59dLCu0LEu7X9vMpEGIWF3leC8/A1Fbd1/v0LPzDpgIuc/9095G/lf
ErcUZpvjYLzEWpmAevFnl/ezBtNDNdeUEbgoDsbulGv8+Zr6EeEdIY1mdxIFegnGffpSNnlIh1DA
ATW1KYA6xvU8ZZjkuWsDvBHhxDj+ReL3hrTXaZUsc0BXR8Ip7+oWkjOgyzLNQPGoFr2UIjGIb9GY
YMUEl73zS20U4xrrMSzaXBX9C4f9/+9V6PrOPOP0tJVU7U4z5BfzY5iQHldljIQYp6y70KT8ODAU
NXQ0DuI2Da+m0warWwnvw4ZG4Gtn93MdvMQq3HQEST+BbD/DpdfTFNTBtQTSfQrnEWRuylFYkhcA
oUkFeIXCLd8xb/rZEES/E5fuL5Vw3w2oz8uND+jng1wuRf9+EmIzGZLavrXKLRy7/TYlyhdSNVAv
A9CKc52IigZZCM6HNFf8jH6aAZacdU3J8AkEQ9XAZjlD6EDU3jARluV9zK4E8jLJLJpz5aTxb1F5
OzVeuwvZuUGrq0Dluwzwu+juif5DlR3HDp5awMtAPM4P+Z+8bsn8qb+ZhWH0zxn7rRoJgDTuBx3J
98GSFzJMEAWbRgN4FyIClhm6A1gc0fWyP+1+EWAp4DhQFBZuoolXw+y1puHzV198bHAbHL8OqT09
TAAvgMrdbEgNmMqRdd38vVdSf06v8faJ2Fx0HnmFT+D1uw1ALEx3jdEKQrIyMsw3NGaXo+PqzODo
Ms614jhsqmlwcEKms1bySjmA5PKTvjSSt3uFNlHLAlTA4P5niWs5gZArY2p53tIva13IcNz9R36O
JRd6e+9b2syGU/Jjs1svVq0v3zKgiVKvyphTjFKEJiJy5ISrT4T/Q2XbYFSu7hmGQYUSfBOwGKDd
/5brOhhkomaXI0G5XbUCSI1CPY7p37GNRhfcFXDLUzTkgLcjsiMXwFXovENfmrBkW2cXMzpQumWR
8jIjjZDUv0J/2SK+/VG/4zOTmzScpf4PWubt5ZgDMVxSmW0A9kW+8rY6H6ATj9oEgfoPKP3MZbPT
MAkNnOlMlIHWHlTHfSpDTlJGrWcS669hlv892mJXepADhtOQZkMNcsmJqX+n/WeilGgU+gERg33D
JNPkFoedSXrPwEd1StRqBhot3aMvDEU4c+HvA6b264+7+ZXhASMHsj7u46DhqglahV/tybZOMrv5
sRvwJc5WV0t0vQH3J3BasxSd81mPqccOTk1FzVmzB7/rSxihOoFSQHkcJNdTfkC/FS1YqS9mXfyB
JiGhR/+9zpIivJWJmxsb+GamJ/uFHQJSKVtQZa7LDjbSr4jYA8KPXfq3AhVe8mmRzC9UrGo1JnBV
hyxRKPxoVxxVDU8DJLayv0nY/jMyXwCovW95AOehdyeLkpuZjL3EofBS84rRH0YFjXTZTGP2TCGm
aP0SQ6yeH/sSG7k+MKIkfbPnrr8M3uBY1e7cI+gVy5DbkaW6gewAnk2UqzgfR2T19XV7RrB4Rbtg
nDrD05kTKRHo2wBskPZuwIvIppcxHO9LHUIitwxL4fjPmN2XOLkMVXqaDCp9ok17BO+VsM9QyL/e
biCXcRYMb4NG6RdJ11pniwREawG2IlbXDSTqy+vVVUFHQTBJeWydHtzdGooGvk9GBRqG7jy0ziOj
Y9wiyOqJT5uSKnu1x1ZFF6XwjD45PsoWjZvdIWFob7gdiDGbMX0I1/zJa7vw06ExoeCf8LopkcL1
EGtAUif/fLZu3RakABbDM3ebI09EObbtKqM6PRuYYIz9WMInbUtwqCnUwTtNDCqnXuDuWPxakXHF
4OmXTMiK8hREq44UctGRQ7A1zGFx/CxK+8T8ipu4fkb+RrCFp8rno3bji9AGBn4NQOxRlfUzV1Xa
KgbsZaIZiZXudmX2AnyVGCyqKgBL5URhHeorU1EMyJ9qr49UtyotXTEZnbPz4o5C6HXrGmgBp2MM
39m9+DXdtPjFdure0XxURbeSIqJOo/vqnTSiPuECsCGSudUHOw/ckJCM43hr8He4Oh8vPszdnbEw
dCoqoM+HBmCoUpY33aJ5094x3w537kxONntjBqh5PJa4w6egAjbh+JHwJVqoxCv7f9IR6MgLtomG
Rdvy8Np/BokoyrRu4pv0Eg6kCSHKsbojWcjs+11jU8Ohwz0C/sFBO4ppJwvvBm1F10rkutjmACTL
yQyuNqG+GzgTnNIOX8jW3iKR3dwvz3eTvcTr/0Z48VSHgokQ1CO1qGbMWtNnmPo+7xLjZCxWvPSW
u69YZAERuyfo0EaNlzVkzBVU8xGGGaWrP3xm4A49crDCktm9Ti+OaWiNWa1phB+SgUlve852kriA
L1F26Ux6hSNjfjqzaHwcGFdCxrxQBIReYrOS/3U1Z96fdB1yvBxU0fz01JepE3CGui+J/4xfkaeo
gtlG8gl5V9E1joYSZR/rB1ZAXN2DfMSk7NoRxglu0GHXLEqnXSCFA6RJRN/mCxJyUUcTHeKuZxVN
z6w4X6hInpBFOxFmbmS6q9eAf9/U+HfqgVuxb6odBtmIBCcei2niz1oOkHcv2fZmbb6OV+kqTwcc
V6WhfstJdwMTHbSv5obcMnWOTQGKuK6t8MhzsqEmkerigfug9yA2R/BTm9rNgu8OBTXqDjPkSTaK
c/pXRJ7w+tCabgQxbaLsHbE3o5qFG/wizv/hvGjhcd8YsbgK4nlNP+QT4uy3TAJJ0RRqtiGEZ1+O
l2MOwAHSUWzGI/js8H2rauX80rsD8lFshP575gihKAaw0w/WzSwaOeFGTuezliTUjPX8MGm7vEwA
vautTYnwB5+XoV2gkSYrcn/LjQ5dFOEfsJaHfY9y1h2szl0ezh5yphe2vypZxm55DNnrb23AHO9L
Qbux2oc/3EE3E6pl779XkmK2Vk3dM+z+c1OjixIMmf7kO0s1k+vtjaYqE1oxbrRJ3mACdfdtlxNM
7qmuiY84WYqwL0ExwIAz7S6x/3HMpfRbE3Az2Emm6TrfEoxCY7fLEjkDtoxgK0YAfn7ixtebYfoH
lX1wRmSerZJH1SUn7zRfOZpmzLZFIWsFBzJnpOOGXapktuEjI5hjAJ2iwbn6Vg2bwaUhNWfbf81i
VO9FJYT46e6gRzcMz+wkUwqqkhRsk5NOeNAIfcuzUgefCWBA84kgOKyuEpv+MsVOOBNSf6it49rZ
tlBfvBg5LsK7/OfpOqh/Nry9WRwOfCM6kh3rgO2gys3QZC3v5F3qVua7N2nKy5UhC9BJdkHVOdv1
+kus27TNrSWuclZEtnFzEbY9lQxsWD1L5oFl9AWYYepYTBtPf3PD3nsq/txZKK2Z3AlDAhFa7WPi
HHxgxSBfBUxxjtWSLphG/wYyc39qxeCr3sOV1//Uoj4G+tc6x31xg7LIaS0lYWFxYbeWjANF+QMP
QxtuUwxLjOwoxzT7WGLWcnqRKs6RX0a37V/u8dGMIhowXnpHvRxy3aRt75SqSd5AEvf7NtZJo9Tz
BS9CBg39rphvHdZLQJrp0AIu+qD64gf4mKWMbOBziQ9ZiuU4d0mIOqeyfoxWu012HdJcA5w5NY/O
fMltJ6iZ3KzxEHaOsoIBTZ1ZmQPUk1WvSFC1uRLEy57DoSB8QWtwL5bDpG5khBI5MhD+zhPChKPM
9UKTMQw2zCkBUBzzU0ytIv0IlEMCmS3w1gBEh7v0tNXRe3AzH22pGeoLtahZAJ4booeqOYlD+eQm
tcoPsVfPIHrW1Y8FPrSsmy2UpcsJVi34SceMul+ZK2MRprz46FZG9xgHsAf7jKAT6Xbk4LaeYhAQ
06ZrxOcaBnvxUXXBbRY/n38V5/cwdM9JBZj3XGk3IgaRlZFHcIrXc4OXeaUv84d6v+RVVsKkgaoY
Zk1nHGwvqp9LQNkPT6Y8f2wV9meaJJY4tBAlNdpfAIBHcX5D/53HvvWPxrYL0HGj2LENUcak40vo
/dsE0bvvIoUfxUAS0t3ihCfHcZJBLnavtegRwnUS10VmebAs3nfG9IMhtphojBZqWRNW8gQiZlD9
Q5PbG7u/PddpPzFcR2dO3c61C5TxsQlrT2zbsnmlf5SdNFoxqaMtSJl/OW3AE0wif8/hLnTut18t
EawDjdAhGpDg3RkymuBwi11L0CHTAmraZFUO7cIMQeHesL2XWHwkTEg7hZNGf7+UmN5IatNunVvg
c7wqrhjuvw+EIqRy1XUHWyuJrFl1HYdoWfU2Oad5hpfFShUGByKG0qBw9jhNj+YFWfmFzGbE9qLh
V9kDlcxbacEk1VCZnZT6AZ9SKTHOc/DgGgMhjYe0v90pEI0rHwRs/ErpFMy6tix8RSmpiEVtEDNY
dL16Dmo/XJ7Pouw1pZqRtm8QfoY6Mn0laO9NbzwUVupcg0e5oKs01TjWVkk6KXGkXYWpf1lUTPcn
jB8wbT1kn5VXJGEG7aJpYVQL2VP/pUdaoFuU7wwFI7Yy039fI5alwjjeBYQZ/CG72HKB2elQEBnG
mJ7WwN3hlbJQA3e8ng9kzlQEnkAgMP3f8B6VMRXDZ1u/YX5HTNzT5ydHLwDDAO/a87z2hD13vM9R
YIb4NwM0WGsWBkm6oHlqqW3mc16du72V+UxHjmNKgTkd75C/sl8xjLBjYCZQ9hDqSkcDUZPLBRHN
9abtX8vb/nyiov98y5AT5wpp+f1Y10vS1qGQzV3IAmZk+YCnK+FN4tGY9CPVMM+txGAJd14sKNQr
Q3jiTG3ayj6zxaVDPQAPux6J8L+h3oo2g9ehQTF0AATRzJSi2STHXtRog389fY/o5CMt1ZVE8rgt
7CBob0phMku4k/Q+SadLDG0pbbSnBjGvbB2JHoVDSvA58Gyhmk8uCklc5FM+5j2RzNFjutJg2dQk
br4OvVxWBpWGwSU1k+h7BbPmAidvGyipeizR4rbl3zq/YDsYrQ8+slIzeqnkrtmpMGmD7vJcGbmL
B2Xl3FooIdtWqGl49LK571DtNt6Y7Y4qsuYQ+CRSh6CTU31wamHjnXu+JrdGUApg3J7A5TbJ5BBl
tAba7Amdh7URg8vRjkqbXpp3EuEli0CCITzYpC05/yeqbuYU1i0T5poA9R/JuMsbEmvsth5mLVd+
qelW+HRQjEfLqQi8W9Qq1JovZCd5ymVj84TvG4e+AwabmCOrtqdK08S2zYAkf5t7m8MSuMH1XY61
SP+ZwdW8JpSegxTOwgBaqyg9qtlz72IdLsr6/GkeNIa9aiozQZZy5T6BQMWpmQP4xIuv9O+M1/hm
TE/UMwdypO92gp0TfQH0SE7ANVCJM8tSDFuLkPfLCok3EHTZcGMcsNwZ/ZM2M9moQhY0vaCF3vwp
jgk7Bj1PxTR1/yW8QkiXXNBY8xan1gkRtO1uFsH8uJ4Yo5TVZQqzuXiD4R48i/irtubxOjOCGMlQ
9NxID+0TnN2EXzS/s5NwfYMNEQmZ999zyjtAlmmRewguTtDLBU5QLth3tEH7/OicDkuXt/hm0fjQ
xAQWTpFkvezBfCVjQbSv4X+F1+S8YAhMV8bnOgengOr3WsSWEUx7Uc0thHApp6WcdiQTJ0zIKu45
yk4G54JX+2zxbpzM+yuWE/ufwmwpILwm0y8m9sZROj9Awv+v/5jN5c66ravAa0GczJLvXp+mVCyq
Y4CDhsG17Ts23uE0RMQ8D3q6CZDT8BgqyVdt0RrawVwym/3EekVy5cOf06p+xIX6ovpBWsoPOjR9
AIFImJXyduxAYKTCI7NlxA6iQWaEc9Ld+1KKtxVqMKdqvCVyaAdrMLNgVlVVh7hmRYqMovq4XHXo
MF60phps4Ud4pmNYdrzvQFdvVQjSXARNKrs0HA2We+ZZhCPaVXIeDTOWmU2Q5Y1buPe3eLjf+WCL
LNjt/XgNmvSO7kxqjQsBtE9EEJx0pWFetFUxbyNf72w1jk8lHndm3GknS2mGbV9aePe0eXbcHISQ
Q7D7tKRjotcOVG7ATJ7WFNHsR6zFIolxGOB8fIqftcMkeI7kA6trxPuYw4fW0Crztfsgo0TWk0as
hUMn315n4DwZChlV7QS4QEgRedCG5EenopHeHQmCqDO/eJGRRgWGahfr9Lwm9wwXH8pKejraBR0B
g4SHP7srZmXs+4m2Wk8yU5+IicMR8eiJG5tMICe9Atb8J5a7s6DjGCz5dKjj1+FrjgimcZA4xPVn
qDe/pOkjcXoPAepHY9jfDBe4mL5iYVuIpyfYSW+9hXQ2NyenXpXerpnDz6VMgEvHY99Nrr+0Zakc
9hDCXDMF3mBifnGda8oVelNTUaN2Ok68/4ROuXSN8OsxO7iA97PWh1w6NGRVLjsp8v+K51jU4ikh
M/bwBGELV5fMJIe4dHGCHcJ2zLzMKiPNFxoE4NNQiSH18MQQNzpWQuAgyVQSJPEM3UwZqubxMwsi
K13DZ7CvIMQRnhtpZUkIX6MQthA2mUdWVq+thqXPxrqhrJKQgRTzSEBd45m9KuQFLONQSGAmZzC8
MXY94DkOMxaPtScudBzUCmrzsRu+PZPvFfX7nc5Z4axsLjzBow/VKBMt71dG2TVIOEJIHFepDPqz
OKeienhU4PHbnq38O+tabknYcvOZcdu0dymxIzeVBvfWTWGVYCh2H9rkrL0NHyLvDGlx0fmUVLz7
kUgctSplra+BhK3Gx0wNtrXtiKJkhqy/1S8O45vf3bxjFUbfr4iYdoWzHaZSGZaRQMtBA9WIlBTz
ED2PUL4PtAAMu+aGu7f5TQ4huSEItvNE5jLRV76KKPhZ7jrWPByHHJjNegI2o66byMAMs/lwc8NJ
ozcYmn5X3RmHBPfWwAhSWaZwqjQyrgJGFHNh3PFyqg1qRI+E4LKdybl64tx/C1rGMtJ3fBlxgK5G
6rHsQpRuEVt5kdTQFtpFR7g+lWE0Ii8nmVKV7CL3NOZzKbSbcOto1yM2dGQTnhNIehNJJYpR+KYZ
bWCK/0Y2wmgtAyg+jG4l/VT45yMafDS7mG0NAVsBCbyucXdrlu/4uShmSrJzPmGRYrLFYOs89DTd
gq7EMG7n0SfWx8KbYIzHh2XpTODXkY2NG+FuNEoGwZwd7bJE0mShB7q+wUfWad1xWmLelzsVga9p
ZSndIDA09RxfFnahC7SFR5JUWo5rLnKo6aTP2IKeLur7Ew84XXLxRZ9/mBS5q64PlKluBky59Wyl
fX0wheArHpXt/ZnCHYh3EOZm0WhrEu4wm5py9TTI6K3jnmL9DCGGZcGESAxp/hOTqyksaOZ9UsBl
JPzm2ETXlq8O+R40woxejLCpX77smE7KkB5muZCqC7hANugnMElF7nu/KYez1D+aZDxAHd8lYYo5
VcSpd7A+VEwo8RF4kv+WuNlwCzvQnlJl+g4ZFSTGCDMQWnbiU5CD20w+cXD4ZsuxGTFvCE6Pzy28
anXKlUUrTy60uauM9fvW6tO4numuzp3BoY1oqjLJjc4ETJn5eB3PD7eraueFaQC8fdvIwNozlp0d
LJu+nih78rJLBNs93QM7hrKRirlpkxAA3HFTzz6JOR6o8tvcPDW9FW/fskR6GbsglTS2qn30cwHY
P5+3prDSniqUz9cD24bx555O5TYWGfoIsd0+AJIxhwNxAeE8P5MtNtZfbbEx5S5KJ1wLN/VcnuL+
7WLnWVNHRU1iq8YtsnCX+avCbP73FpgWv3MkZVlo4fZafonnl2kPM4ETOcP+zReCNlawBN5hRV0v
gnvk10FUf25PRWccEYZIK2Xe/qDZbhGybIIMM7rK2+BX6p0D9348G3yF2cCefORz+VlGDMpNDsN/
yWeMY/1TkAMlyfOmzhEWnixRpSyyhjh9lH86kfINoAjzNB5pKREvXhsjlUTHYvO0IyVaUflClTYc
wp8mCV+y8ey4FIqu9Q20SkoG5eBKsBCS77PlGfXTVwS186fgxql7RNRDquTC6DKFupN8lgSWuUro
EPlgl87xTPBj4Xpxeab5eKbmw9ne3eoSTJZQ2fNKYymYTaCc81xIt18u03CQTuuu3BWOr5fd0eFH
AZi77L/J/uTPSMIAtxyVDbxv532WjbXMufhGS13JCmMCiFOBFsShBQS/2ZebMq2OvtzEO28OVLFg
BfgtVd9+f28U8VVz2XqDSOZtACeIsRh/EzJL+6vL7WRtK+iazVhi9cg8ibteEvOlPnTQ5Ouc42zI
UhDvW5TjYdIBabUno4E4R8+oTmL2TU2CNEgENNf74oK21ot/AzbUfDdcYAzLKoFQPLtDpvVwrYne
zc2NIqr94eNx5nfYQXAhYDloJUXfrhbEiok5fk5lW/aVCcbw5NzyB/I3o/Qp2w0HMzduw7U6r9ll
kmTooLaOyssO7BeKgtkzeYaFywWU3scjZo0SbXub2sj0XMAUZRUOJ3rKgAmLjOJt7ObS0xzoZiII
nT8RZzH29otP8pE9tBesM695Jwj7YeOR+YuRv/WwQxFYTDOzbjTfsa1IgyORUJB/exhW5btlwtuB
h8Fi8a4ekRxPy/mFWP8AHGQ+L95xRC0yxIs7PRKB0HPbA2epLC9c2Y9QSOu+iqQRGm23nIHx8X3K
qQawRTLjJXIvnUZSapBHBQfN22m7tF32psN2WzTVC7CYH1fG3h3UE5yFsLAOY9dG7JZCUDM0fFbn
2SSSSJ9eabeUdmg6B/9SessuhwaSVijkLbiirhduzOoqJc5hcJvTdhWvCHlap1FMT8beXA1VN23J
LtzxKyCNf64i7br7MbopUDyrIo96SKkCrLydHWHQ6j347Bc7r3jcL0H5897YzZ4g1Zla/VVfIAZo
L0Q5nL+bTdCQA31qrWyVIHehR/BlP/oVz8iebEy+cm52SvqLmjj43i/wR9SvEdbIOfJk8GpavE3b
Ebg8G4Mi6//w0/2bd947RCrNP138KkmPvnKqb78gDXBegyvY4LpxwWUh4YxUNoohVEwACd0ypy2P
PILgmfxvbXDO9uA2ExX/05zMu9lce8u0okFp93NYgHQFloE+NlMSaf8zdalez+BNLlO4u7NDnv/6
qq+e0psqvSRzIUH7LlG0c2alzhJWlxDMNQVPCoo2xoYTwMwYyz2lW8WPZCl7jc3wmkKykT5KMvsq
Bv9DcYVBui2YNUiBn4jGkr3bk46j0r5iSTfO6e9r5slglEdI/f0y0Chvahy/8TOdsIFv+VtDHQrg
3ySVEZZWn5I5f+TmJL70Mn2lJrA7WPK89Qu91iqSTYnUl9EySw4rbdDWOSR6jtooAG5IfM6qB2K3
xwVYNXY85zqYgL6mvlzBYj45+zqXhB9WIfj9A5EZ1Lbt63KeQUCooCvgN/SQen1qX6pkAZ/WUZIk
I3Cg2+n9X7wQSt9+BotbVMOr4ng6ofwqfwaoUPRageHxl6YF0MJhkXKNFpE54hXoYhotudniY18d
nYFmckC+s/7hmYbxwFG51BdyC2ZDPGP68QZICbjwb+pyM8X/xkF5qdxF0A9Ka1CGOwNvnhoTJLEL
dSERO3rj9G/TZC+GAoCZL2yJ6IHJ7tDg3sDqtV6lnD4oS1fnMffSY8HEMxSAR/EZhRnZGDt2vPv3
fylRdqcEl2x1kUG/DR0BxCbjxWwk0aVJ0i+tsSfQqdB8w18oHrCLo0KY/P1EGSqrrl7aT72zBwjn
ZdgWAdT/RtcOewFnyVEjzrf73W3ie197lMjbT5x0YuNUSSy7FgC+TAAKuofEIPglAUT9dxxbIYCk
ps8KEpiyGPe9khczlTM1OFWL/eF72jiOSQxXVGZ1XRuap61ZAo8ysHrKyx3hsilkZPlztvDiBfgZ
LZe3jmXOzodEgl1y232WXgzx+bxcMW6+e3lo9E32V5BvZwwpR2B6KRYTuBSG5WZPyuts/NNMosuT
xAJqrbUQBV99/H6DZJRE0hOfkEdk+DfnTVtQV1AcdBiyCHRhbhhYb/pp4S6MVqdNU+hedlmjP8ol
brQnP+SK1Um13elHCKN6hwspm5LWMyGunVdFEaiVMLukUXB9YzKvFil8zJqFLgURBU5U36JftWLL
yWMrjWdDt/h42jkih4VDP4BnEg46kdXX5ngIA/XgHLxNqCeDCTeM6n0FBZ+n3mrxWd4Aizvd4bK3
GuH/MSoHmU6jKiEQujgOLzs/NR06sk5+LbUxfZ1xZIqWhat2puW65sO7dcSPogO0OC/M6Za1LS4C
SXMC9Fo5J2BVHtipEv+JAXQvSOsgEUNWWS9eXVtzK6t/opd75NYFpf3Gr7rbIwxEU4Z5xrE+IAT4
kaeRsHoLvVWvP+TwB+SKeBTcZdkUHkyjgoiqxuEoFdD8DS21YmddftIfS4RUgALmTJKJSjn3+qOz
BJ12vToUsbz5vPyTLjWChc8biE+tTxuCcar2NdBFocYKRT171A6tugK1XA23rTDGru8D6yclNgEZ
DdbCC+N7COitsfCsN5FySAJwe5je3aBtJjmP5a3vHJg6Jraf7cP/hTnXB7r5xKJtOULUYokAEbqI
Xk5XTXXZwsJxFCayCyqMY/eQgZM0vwVWAPEFaldHmT7r5iIipHqnZuRP9gsKyIve+3bfLBUROeGn
VXu/VBQ1CgLPaG16uR9qoOhtEwblDUkmVGcsjj67rhHKnTE1hKbiJAozzH89P8nedT7lHluM8YaK
mesTQO+82Cps/Hb9aSw0BZKgfL9GvAr3Z5W84IgwxUfK2SQ8a4VHDqjqFXNvVp+maA71FW8vEh2c
DulXu2Gnrm6BW0f/+S3ePRaviZL9Y7bDuKdnSNkpnEq5E5l9owieAkh9o33XYAwnG8cEi+9CIO46
MaykIV3G9o28UTWIncEbbzxliHHg3LAU0/y7TIrBCvo9bCvt+zYgMl//uYgoi1H6LzCjJwqMPMCy
sIThhRalNZgbHozId0aHA7aFW5yI0JOe2qa/dF+4ULzxKVXGBaQHl2WJOFZxOVS+naym5pZTB/+T
4h7HdtoBkIeB+4YTbgGubjkZvqoQ4cR3mCP5hi13Q42z5fYIp9AqOhBWGFh9LqbP+DY8tq/hqiSI
XZ6X0b5NRKlYF1DeSt5ZPoJ3yL3BsvuiaTKYAZDFY1RPZD+WkwwNK6ETMnVQaL4QBc2/2ln2BuWs
eBlbKmRMU7pvn28gqVvzOrp3ui4qO+CcZ/Kaqs/LN9SNpTph3Vyo1zzsm1Aq6S1OTxAxlk/tGTkW
nPHY38RX5DNbnDnERpFa2KTZkZKNxpesHO4DXhRGbGR64nzfXVHt2/8GYFZdlibjCy6+4rFxdp3l
yQDl8nSQUmKbgnLboI5ruQnZXfLJ2PSct3B44zC330NR0yIzqDPch2bOfG6D47glIDgLzp2dYpot
nY0oW+s2zat0S8aDQLaGuRYokXFfENlg5w2BOxpJ11C2e7Dq9kWCavqfNcIo7WcmBst/a24tgXmi
PXb3VDoRJJXehqETquRPgt+SVAdzD+g2FWUshR/mYKDClVpg10bqbs8G9t+3cmRp+eC20Ley1LAE
fmP3L6oZ7JVNeWeLUbLBT94vvQuxFCP6Wftb6hLFCspzq8coS378+5Pr2aDvvW7hatdaO5fsLrvd
aSUfMKT4Ku7qvQybyE3VM8ttFXkkOXeHGkqP5yo4UWKtkQ3QkJmN+414Q30hkdjpY9rop29Bn9b8
w7H2/mOLF5Qbb/2esJwS3W1Gufc74N0TmRAFNENycV6sqtkg1u01m3Kzxu9pvIsIpraMJ1slRjdV
MyBaoLiV0vTrRjFOVdJymimcdxLl2V/k2BChFINqb+QUVsyY6JUsVc1AYkvmoDA9XZDXzB+eZUL/
vfiQcj2nxxPyxV0B6aFyc/TzcTvUw/pAuU4YXQgEkK8N3nDI/U/6hLr8eseRhWDy2fNXXs35lh1I
cusnYt7H8faon8sDvdmwFIubhbQxRDbRfPBU69//Qu+2qalLyNYTv+jtG4W5R4gNl1qI5TA7Qq5c
GVuMyhIhvDTuTCiQ2qSXxKy16kDXwWD82k0VhCRIelJyiY7ujntWQC9REmAywBmF7XzLyha8t161
euV2b7ZIjRcG3UsDrzz3M3+l+zOsao8Feg/QOuFQAE+3qfvcgKPl++LQmWfJ/pOpRebXKjnOY+3T
pAWsEHsqCoU+E6XcOWBqXPDfo08Lb3on0QETBBeZjCJX5kP4SCFvH6yW9wo6KRuOAP+0O2Q5TFWs
8/Tnh2VRmFaBNw0pi+WpYDc/ocEiHZ//6NyIqpIGuQHInKiUQlT7dmKqco96oODwMpn7Tk8WjQgP
1YvOcd81m5hugvg++w/oxPNswyPP4jLJFnMPJVcs9lzism79/A0PGYbNcoglLVAeQBYXbWNlPv26
54gQ5PBWFN0e+fh5UnSKOc/wv3zJhfYP21Zr8zViPnYb5pxy0mhbNpXuAVZnGP4Ej1n86/kxZXOh
++uIZyQ6D4vD03CgY0aLE7fsGPlyUO3Y1KW7l685riL05mJOFJ6kXGBAh7BfhR55tkEBuQp1AiIP
E0ahWQRG9KsIBv3DyX+eXCD8znJWNBgUh+9p99lz36Hg/l7vZtZdPmE+Wk/15kuhtM1kh8X/sCdq
yEG3HF1vfaXsyXSml9MyzBD6esmYCA4aI7O3PsHRKixZmGEH3kO0+k4mDJY2iWGBf4YBZrlH5aMD
XzSD84CbvJi+Y/Z2FJq1WU2n56jZgWEz5baf8Nau1SNzX0XwiZtCFHVjd7VSp3NBiB1GjxH++oeg
B4Isyh+jJNWqtLwWyvGpN872FLcJYPyueO1RvZymoq3yBDqawTsKKvFF2UOO3DlS5Zoh/7r60YuM
/3+xBM/wDMR9zLVHQXWKq2omQmxgbRUdPtp5EgdotnfTgfVFVZATgRfgztEjAQfcWkzT+IkJyV48
8C5YJpitvt2wJs4epGMjPg/MN3aHoQ2gk31ATZFk8AF1wFCjT/ateN5CWXrLoAwL5naMV9b0TKUG
C7/GDhZxiA9XPkqE8fMIWGtoo9nMoe063ABbBAs7E8JtscNCm97Z/fN9hZ5F4yQIEusH5VYdWGCu
RBH9zH0RfhpNmwJggxKW5kSOcrvAxVSW1pfNhKVuQXowgXxUnXnUSYChqRlyJk0ldhxDwkNhUWAp
XCt7UssP5JfM5YCNyj2HE5BHDBFutOrTDtUDMMS+9FIDN0Mv5B1nDU15REqwvasJElSYaEKaJ1jE
H3zgIQh2EpVSh3Y7qlfvcn8nvPZ7XIYR124ta56X8fkMP4BzYUR+ZxbvS9lE5QmH3G84Pe8nOZKA
fvhyc72TKn8eVU5pGNQj/YnKVCqiMpauJOgyPoM65P7hwedEHi9n1KhYBC5h3kISCb225AaM/W7u
g2SuW/vWEq/0OW9DM369pe3S36LBFioZEjmqa0Je6KUeRTlII+IRTaVmG+gCyMROlzbn6mxexOGf
sKxArksQsXN6WmgLzNBTI+gm+w4pFX35R9AsPefWHq97smVYetc+P8fnGRYn6qleJG3Ex22oiio3
BacRP3KH6+c/UjnIvWSWjKjDng36a3LkoRQRVVP0H+WxTpFY6kPUY5vCnBVc9t2BDeV4caCOamik
QN5WY9j/ibygUwwMgq8BFjFmPXMobUAQ++AF8c2g48IDmi1VNWsG1e4g0TsryN4KkRRPL2LTFyTG
qr8WmB3/H/orLwSj9pe3WhLR0GtJR0PS7yqsJycX572IxK5Gz9vrpjjVyhiPSf8RSCTuAUTPYI2s
lT+bBifKDgX/TncpXlFo3Ng8AozbakhDCjnoq83OS6DHo+9Ozmm7QhGfsvilPakiGN34+XGOIeRR
qkWntDoJV8k+sE8/iBFjCUhEkzJWfHl4yCie+dYFTdWCrNZolXm7YflLIKEac0plg4Mk7EB31ugY
5ZWE3tou3CQFDc3zht0I9mLqslxp7LsdRA1423fuljkxqbmVI5Q03/y9nML6Kg3TwsiNIMgOK5ek
YomBbPVnrGPnUSAZlMtHKHbWg64mPTwrBcg47HZWePqlkRbFf0E1peThPpn/WAEzqPKF8mbJ6BoX
nlhExBKoM7DxwW/3wdWHKHs/5SAxg2pNL562OgJdxCR2tFWG+cHvEx7NOqHHuklvWKVlHxpZJHFT
UEsAyPYvmPazDjfjc/gnOeZknPFMiR3b7n+LU3mjWB3ALSjzSvglXWPrF+DL95mWT5H17BOier4x
TEljCNW07uLIa7iEpNx5KEOhinXolfLqjxYx2RpsBhuAgAMhJ0RMOfqe9BY14HlEigMtOTGKb2T8
f9FD/8bqJ7tFwLpdpB9WSUyFxj3pcPePfna2os40nRR3h5Q+lduydET6P2ab6pH6+P5UNCQAKcTN
yw5GsYoqt5hIvHQt7A/H01hEu0mTHMcK+IkXjyCZw8QKllX3TMUO/9hzlLLESG2QhKPo0jSzTgYN
j/7319Jew+SfTARXjB8wQMXD8FsFilEMhZbNuR9v7W4P/4l3pie+pgXi17mjUr1ROHdSkyEKEEev
Y5r/D6LX58BYhnC8UoX5Mb7eQxSe/lv/pqOL4OK3zm71vq/oS65vMXbm4DMz15Lee6HHTiwaD9CM
KeVHTqQT7d4mWdH615TVE462Y5LP1JGAy/B3JFKM1k4gW7dDCpcX0muzSg/LVnEmHqViLtJHbgeR
a0K5LfKv/Nn+9pjh2JORsbJ3POzfpl6rPQjaQeuJmsqhlWFmNh38pUizWRDiZtLFwe+hAIbZEE+c
siaoxdUbXc3iAe3P2VTsaj0+BcnuKxuJuvb1FFRRAJlPAHjHWB7/L6HNs+SCL9KbzgDzPcyuqBF/
GSuOYxpC+A91VIQ2WSci64HOc/kTMFDMJrtZj8XDUdh4QDiCU9anz8oLIfAd8ivrShFVbUid6BEf
wkwV4r9B9JMTuibgq+Un053O0sjiTAQDvQwXoepR6HX63mFJFdTsxI7SWS4hA4F+ElLPEKXmI4XX
G3d1Ce3gpwlclb+vOXeeY4CcvtjlMJ7WJTbawQW5Q0Ogzg4+oPxxjW5/NvcO22JszfVoVwlk9UX5
IIFhVVpVRVCZCsuf1ES5iWisuwJjPoSxiBV8g+uJ3RvPnX7fBu8esuw4v/AKxhNDgs+rfFw8Jcap
QtdL4Ymj6jxvebiXVDcsrvnMWZLFItXP35C7+oyS8dSIQxu2KkGk6uYyfEQ1t9cjG7HjDhgoDGTN
Bvp6msuTO12AVNlQzpPgC3dYJReJkXe3rPTw05LL8gXKFe1HvDHRCx0V4LJ9BTGoJ404uMmGOeu8
nWkxgWeta/JOi69KkNtO7VL8OnPmq/ceiIWEOaw/zFSA0vEOfHQqfpmAqezh3SoR6Sr5cGs8okOK
ypjr/56F6DO5KQngJrcChZQCmtSmMEoZHylBI3CoFamhhT8vfakq/An2U3gJ+yFU9DvlXr7vbWbl
Br3XHDS0RQf2vhZ/sj79FXvMLUYB45NAYMTEORCfAVuRsxiA6SPfGwp4lwwJnSmjT5BHehV8auTb
7DvJ+X842VkJXxQix21CLI48eG0oLRkQD3JLz7vQMFJFcAjSqWMGuuLgbz6dviBOHgtK/sHLmqcy
P8XUkJJ2fPTzSP/mGiNzeocDXxAkBTUU5YBAVevfOV25N6mwza16I02+rIon1/JSgn6OyHcHyYYR
qCGfJxcVZP/pUg1UGqvUXifxPFjQSYZFrni7Z7rjlP6IYAWfXjwYyM2yJ0ZeH4aP6vfqbZsESRCP
NCK09rH03lwsYLG05Ri+dVQpz/c3yXh86zP1jFiGN3bgdRIav0+++nmtq+4D8jJW/U8mv2wK9Y3p
EOW2YRDAeGrulR/I7IXZeIwaWVU7vQKLVlYA/X1gKvYfMjXzodUR17jt9BGgFCI1c9q29Y3eV0s9
kGnA9IOsyTlcl5lNstXQMfvTqo8iEcoWv/dWSHtDU3Z+TxVLyChSpYI9s/ti9QeLyJdOT716o2xW
sCakwlszmp5HTM+nncw1UbDH+T74Z8IXldHYlIoCw609KXVzA3wS9QKTJqRdY5FEUxX5n4Bbt4CS
e2AquT1ihoOfk/X25/ZUkmBB8pEOjKZM1KPdXCi6c7xdg+Nb47E2jG20MPdoG+zOnhx8jyjybVh3
/WA0K3f8809qMIVkjnzi8+XsmHwiXD0cWfk8oyHUiPZ+/knoGEx5e3teaU/Epne0G31SLw4ho5iw
fPFOrRV/jQTEnBwAKQnWtZmfeBQTYTb70Cjm5d7KM8ouFjIyEixEUE7zR/n3bCQOH40HnT4jVqLK
pAGeoHqKP+eIMgEoTsR2PPtJGVrf5IF1sqoBlWUkBAtuSx4D/q4XTaORN7u2mKJNfAoQHDfhnTgB
UCa0rK4HWnLWe4vedgrpbm02aroqXZbmjrTKZavmLb+pkpLFGOWXlmCbLF98ZmIVbC0Xee6XmpCb
LSoQOJ+Q40fCTTkvcCFKrqxM2YOJPQ3jGQ2NLf1h2HeLN4Kai625p29MnhMVNj9Pcr2tDB2lN3Y/
fQVrE+MsVxdOMGYsrgmgNir5yG/Z6jKOtTEmIDUrKXQJ60NhfRRJcL5uzAz37qWOIZUGMmT3b9Bm
10oQNA9UfC610D1NHb6iXuTXfQ/lTxrIjMgYCyR6j60J5bsySCh4wKhNAkpy56ja9rpHGNw1qK7U
4sceCabz8j4BHgrvhZkPuYKfaETWwCWxULGZX3USo5BSGmlXeoxC/SpeIt5nXeLS18d+SlU4Dwd5
2MXwHProG1YNUeB03fKNN3PK/kSXbuHyRBmmklDTY85o02vmpHR4LP2xzmFDaP12xUSGlafD84xU
Cg1IGHiv3ap6Q/J8xE2opxfrs28ztwjfigDOL2oaYCMsjBJqIKNfbVvS5WY8VstsQQyxJ3hhUDYN
TYAScob3n9mv2PTwuXyFZ0F5RpybC9SjdRA5X9lSJxIUIYGv1gP/F/7aRAvID//mIqUgzOlJZyEW
tyYA3kKtP1Wr6fA8LqUVw50nAis4FvT8dFsiRzrpz0vlrJn+Oxhh7TLTAksa0YY6jjmqzNMCXxrL
zeH+kJ/sjSLVDZgGmx8clb2aMIHvv2f3EABEIHFGqiW5VSzv0RrFYttoZ864cQOa/eGFOOI2c4fm
MBuEtKrL4rf2yXBfUnFE6rpIG8p2jJq21UpeeK9iGOOmoH5N++YpxxlpAvOwSHxbrDKqJsK80c0c
wHRfSmK34mLp0ch5C3Mt31RdpUrr1tiTT54vSyJRNJRpLTDdiFD/pKFX5XcAY/QJgHxaCJDEOXJv
KT8tQWDSEmQDSVPeTfHoJ8HTMJYzx23sBvp8/GGD1gYt1s3y76tZE5+ettWAklZx0MQajSJom0th
NQEUyTXLhtpGu6BnEmZGHJVJStR05EHwzbTBw3SzF4kG0pNiSkDkXdaU47AYmw4Q7aM7c4x0kpyo
C2cn12nrHQQSEzIAlRshE4khGn6vdMUhFKWcUaFYJNs2syHULnuYmELpawfI/KOHQcMHGVSL7yXK
9WFAy+uPU50se+1FwDxLJZiw4UBHO2kzguTIVkkBlzglZiO8144lLF3NLO7W05azKcr9Ou8MfPgS
nzhDdWTpBjNgzPoqQQwT8t9y0UaA3LPZACZHGYegecqkgOy6Cndq73v4jz9ukh2CJl5yAimPOQ+s
38LI2WtsM/7BHnJVOiQ9Y5uAaD9C6O2YpQi5VKy1GAGco+HCPZHUtmA1HlB7vKhBZz1YW65uZdKf
/tYGf62OPUyDmZmyeu/lD5mexTcVOEAB6+mMGI896Nst54LgF7b+FkXGtpwDC1Sfj7YSesQLKDW3
l7v5mskfFexK9k6wgCYBLKaWtRcgfrZ2QJP/cLQHTCn8lc4xsTyi4V92sLnGOoQkTT+iPkV0a/AN
ME/bmxTMLwo/gcnUcTmQHcrjWp9JFU3xps9twTSzau4xFVoyf81wt2UKvq4PxgEIrGA2SrAxl4Jx
jBVLroEHB2mElMzjEw6ljoUKS17pj1LV6G2N6jjoetZ/YGnRUsG8/QEF03tAMSH8tBIesGgEyeDi
aHm6MDnOiPsU1jmJqqnyYTs8Z/V8D0eVNPdsSQDBE4jC4y9SGnIAuoqrxO6H66Lf1U0FicM/AFj8
c5RKBrZyRm33aKq+bvEW31Nsrk1kp+PJ3bHEiDGifTHeepPek3PZ2ZWSXws7jcSyFeCSGCo+YHPG
9sb8FXsGaOALvPM2mYraz2HP6Q6D50nigunX9Ia6ywL/ORkjK6+YoOGMfXsK2LHXUM0c3305SL9X
01DTGiQsuXGXJubHgAZ15ZLeTlljfEaOj1Qxpq9dXvlOWnzHmQ4FnlfuGOaLL/ING8lzLlR7Xlvx
Jk69hCGsCwAl5kpqwMrCP5VrrNBR4Wasss55RNUvn9yw/7HO4pTF7MScnbfBHwjbOI81Ageba4rX
bBSE3cLL9bHTFhROKnHZuH71PkMBkyn0yrVo75M6MfiKGFJdNZlNVTwp2GLE6eIOXEPCXnfVsYP3
E723Woft2+PEKKFdpZ6YlH/10l81dSnMA4K9P7oV1+DEpN84FwcCgmiHM5NzdSkbyaBdmpAvM/w2
C/F1xRUCbRb3li41cqiB5AhiRygMlCiTiGGYiH78I5G8C251pvjgqPV6LMaDdNqHgw7LkN8R66M2
OPOU/UJUkG7VOfReiluoKil4mIwjdbiS+vqn3ed8FM8PsQfuHPEKeZY+yEaGnjqH0JIcy0KRPK2e
XggjfMmy0VuoeP+5mSqJQ2NCKFfn232ZZDn8AJfQPZqzwjiXp1JldFwK/LjdybVXmZ926LJoNS1n
hZVA4qT+KPzCN9Gc83Jutb0sCgZO4cdhc7N33Dv1Iq/5pGQsyed8SgWbSeRqXYzsprVLn2lcGAPf
W/VcWhKnkbOxnbUVvltcWudNV9DHlY/07IIujuL56LVqX8JBD3b2uvcJlRHxkiVMMdeKosdB/Dd7
ECCzhCGLLHajn2xDOp4fcNgimPEvi8iCGRDYTml2HjvdQR9EzO63SXg6a/kVXjJdhf+M429HxhdT
aE2wHiMO0isOx9v0pn6x8nb41nwyL2wdekgq3p8C2OZssqK4mfCa1B+he3HHAZnn+jCh+zi88BOm
Dlwroot+VQA8LpxG8spVVPow4oBi2RT/3P0c9c6nAQeNQA0Y45mrRWvSasDZ2820RdgPYwU66FHt
kNAaOW7EQmYmvWc9nsxNGsxpe7qr/xSF8p5o3niDWv+ezuTJ/8GDk3ZdhnxNZ7GhqgCb0eyBpC2B
HhSahl1IQCfFs2QV4w8xEayPO5JZ1Et2INeJKEvZO+ZAYQgKOWoxuu7RmAjtWMtB2C921HW5qsVQ
PmrHY7j4TK/OhIRJPFygpafEn5e/zO4sEPMwdpBaqBD2WbsjtPI0QEGbrvQUS6tfxbDNHcN6F7RQ
yqsOtuAK7HXHtXG6kOXgdcZv2bqgeo5Jt8P7jR1nya/mJVI8aSV9ut+sUbth5DD1spCip7qKHjhW
x9+FO6eBsJaL5a2hCeKVHXHKDhTMQPe6RSYUHLI9hYQ34SZLV1FczS+786xSaqzQ/fJL/qTdqhPt
aLhW4Czt9Z1A3teDEGtfwauf9ChsJUQLzkm3XuCV4jVe19hFD9DRhp3xqsTeT5rEgkLkOZhbVtfj
qDrIwXdqcUqblTg64bTpFPbcLBbB0PY5NPMgrVFA8zCk7uZua5ES+x9B2DeWYLCHK3S2nqDsD4sN
SCUXraE/mU1yVHpp55YUffLv5an/bwI+/EotV3O9p5D79YzHdjTqkdb4irjMgwCQlX3538VBObRo
ffLeATQBMUqKTU0DrGM9dLln4qJ6iPSP9KXdOnsoWNQSpgBoKQ/kEmTFpza0lPIGcCLPVEE38Kro
BZ1xSsgytKjHeVzwqHxCDjmsh4m45n3MKavn+X4wqRYUuV5Zb/j55oXrOnYERpxLAyFW2diP3EdB
kuD7ypF1lsBQBcXypB9g6eDxhWwD26jAI3E8INZ/JkVPY6FDyxPVzoIvWry5sMGZBvSkyhxiIit7
UvSfmzr/ttR7Emz/AQrlg8XS23JA8w3yQ/eC7JaTfzdDSB/WfbWJNZDxQ7SmR0mfRPvaKAeCeNxT
r6zPCzulC1KGg+dzYj/oTDbcFcWZmARNDm02QdJDeVDdlXr8wMCkpAkpJ4zmY5/wzLRnxbMgoADD
FzfVowlLhuLYClpFT1LbMeD7CWxPbtrcKxcHZyAPgX/o9xwN2EoS/8q+tcmsRle47Yei7ksDsc1E
oV+ohZlzF9LoiLEjm9WI/deDSDvNYKA8rs3RThyNZQfrrQilgpfUQnOYILfqk/6vzTgB9Dm0Nzs3
FVVHMfS7Nb3u0SFofJeqT4nIRxrIJpHVqUPtJUmN9MEtyzlPCZdb/O0EPj9v4V7TCmTB/yzIfxyF
r/knZ5Rqb5MIOJHBDyka2OX2heE2koGCbfcHm9usRWJ2ROfBCyq6q8d5XJjy3wbsmjN+ORYfuv0p
BPjx2FEGWq8iRltg/SO3m//lK3mzFluueMeATJqlqOVEDnI2z3uJH3GRqB93PbHyIvWP/cPfEAXZ
b1W0N3dcLPDEXP/oeYu//YHU1MamenlAxlBwSXeeJxKux9VNjptYhTrSby2BXasUVoZFBCclwBA2
KyU1q3zPIfw8i1Bhmirp7C/d+RbmxKnHJh/O4NtX6PFO4UOsi1G5AFORqfd9VgzazJKyduRjd0QM
0+qyEErXFwiMyRcfuR4Pl8O6nJwh2XrHFUHQfBQk0YqOdB6MUYhFWUdlvCG0To0jXuso4WpN33+s
Igy7emH/KQiV+mhU3oiJBsktRMffQH69yJwW4Us9mTtyPrdpevzSiGnIW7ibaLJI7QlWJ8QZ7YC6
vcfa66cRqZ3Pmrk4S7t3uaF//4uyTg6hk4von6hJrOImJlXa2L6UtOxfu2nTALNgSimUe1RIwGnh
fjz/cdQ3IQrngm+oBeZfQzDaKLzAllo27biu2Vvc6V0j+hOrF2/LdDmx3B7bk8Eq6UiupaiV3lTd
Ge9lCJRTyVXw/mwg8/L5mwkDwW0z4olbhyPSnVuWhlVNYfTeAqC/kmehcoCzySH4g5wwEwHIUpGH
oiLdzO1iEg+4DFboVGHkjcOkiu43CV++dYsLEa8+IjnVfbbwqz2UYcImUSN8Yy0hA8CXjM1kkNxN
W7dQYPRaPLIeaTgbT9okjlET0XyoqsfyHbzg5EIwyaJQK/I94qnCScwfQM4N2GDSeDV4KMN8FGGc
0bRKpFPGJwQFk6OJw+pQbC/PI78iCZcUk31NeQxpxPFcnxkAAYBjn5S+CKcvgnAfT9rtBQ7zhn+w
su7hxKqVtcTSb4Kny326iEvtzOpK0F0qEOS0ko9B7lTpcDL0uXGhytGMGpTQ5FbLwf5bckQjlrqp
6JQTrSJxJo1lwGxPg9h0IY0NNedh5xXvgreo7BhS9kAZHWsSRIE0L5YT8ugaWtpOqnQFceClencd
ampXgymra5CxcbIPPYt+1RzYajApHTqDYCDiWuV0zA/sZJHlg6ExZ3H09LAnEQbGJwPAdhv8lz3k
wp9jdJmQlgmtBZLtscYa/u1UTjlGdTc9Bd1hBcrazGjuxuHmobGU1p8GaoBq9uhItzW7sZvJxY6W
37knvjMwekz975qL4tU+rH+OZpxz2S5sfTRObrbS4FoRnrEojmSD363HtJpoxD6m4M8EdePDuOZL
cX7FHQGudMXSo31MVlk4G4qsY1T5R0tHuGh6m13zqB/Ayj+worwiVhb7UvZbWk7M+4cZxxNZ8aXT
2TOcJDXVR6sPkkoT3v00ocLBr8cQSNAcBiWUxKC/aBQ+gzMrpES8/T3rdPsFHrPtQ7xhBWsmMw60
FZzQhFAIzUhYC7THvo15QqU3QA87Q2LuMcCG5wlQ2plifKic9W4BOiNopJ5/JUs8/yn7gcALm75N
4m3jXxb39JGfkqn2+zIHxP5L/hCrO2fQT3IqVIy9DLFs1+CqnZnRUIDkeiFsS25wLi0BaHnpdbaU
goDj+bzIONUr294PU/eHkl0ycTzGrRhs34Q2SDoObM9jS/GcxotcbLRpxnkW1sWqglCUtdi+g6ar
vV1BJZeq93eBm6LZJgj8thO00xS+QsKwUEGTA3DjDxoBc+k9ocPbdr1LZDhfSSprX3N/jneQR7po
f7nIc8vUnlv26c3FXl+Gi0r7NeKTst/E6BC9hV5+YZKnXQBX9xjBroqgsjnplJJR2id+piTpt9UP
00uBUwtJYxK/4qMhBpxHwVF+XZwAFx+h6aCgJHsQoBjzz9/qaFD2/y1Ih0LMMBADEBSeWis6yh2H
NCTg6Ywy8+KAEuUmr8l7ZcAHw08pr2/24vJbvw9QwnAcTQfLpfuBz0A43sCenWV9ZBY8/fLCTzJC
Sdxj1TLLsFNA6f/2xJL3ni2Dl8NnBe2yKszjiPxOWlBA/JvLN6ZEHZxSkpV8I50DpCHUiPaA69bi
YWoQFV1epah7MjrxLOVwuum9gbLWjrFiCQ9J+OT8Zl/qKKOzVYp6Qe/6AmNbpyXZYKykqW/O7c5m
Tl4OjXKEjgoaCoqPqqdn+lCQtYMkdir3dGQMAfb2bHOBhFwGhfBltaw4l1LuCFcygBiiUFMDQW2A
Q2R92F6tmTnyTxqSsVHgm2kJfhAM/WdS7ykEoGaTl7xeaceBvrCNI//yjJoh+RylF1QhDw1rkP1f
kqq2o2qNCws2ILeCNhg4uxM35uHjJr9dTvnyTadilZUe1z87EuHRs5uwLeIomtRCzSF29KgEQBJo
AdV1gU2PinqdAVtRiSpQzshzNWvgZ8JtddNbeHsYMMFvZC9AryowiaDWtGMWgODRflq20xJFfBnX
FhFt7uuDgXTnMojr/0jUUbxIwdio4Md8+6pnaHMbH8a23Mqkgt525X21NWGZqhh4AxGO/8Ec+OFk
VXNr1JELkTsiVgRDV+xOVaRUpm+OctbudgRnWPrE5dPIgZ1HA5+poKC2m4yj7z1tAL6afg012tfP
dX0UapW5DMKcaXgL+kewrkNAzxEo5ONV4Aa1ToHU7IAgCCk2Ixzrxr4X7bwEGuqf0lkbWSpweABS
zF6pY58JyRzkXALcoodJioPbM6MOViXXr3/szEXKeoq1gbEnxdv8HQ/vFBSAROsCCaqLKAz5RHOX
4nZtrp1N4s5zLFhCFEGUOOeczKVs9LTQnENJpJEX7RVdV6LACzlv+ZVhGrkbKtSh6bRwlMIDwEnV
pV4N12Uq58UKlwtd88PAIBBSVabMMMuhvFY2EBY1Zg8nY/HnRuthqM5zTPiVAtNjGcI2/mr71En6
F+EqUsoWIG7yerd+3FFzcl1NJP0Ppr1cvE9QGSBK09KPXwXIcMjqpOND4xEGjZR8L6uJCp3P+JhX
sbHN+g5mrFYHDYFaCLTXgurwrYzERhzM8Y+YME6+qIG0h10ZjmAxvYGybenvOMMhTJm2R8TJyr5r
mc0rlYgLNYx3GkumJQaoJlvml6OI/aMmlSLrNprbKeUat07kY0rfba8J+pq/4QvI+5ekDbkCb9CS
y1RbNB0ACF54pRdFJ3Ojr8ABaL4Y6KZIZzvpjtErjBpPsN5NKt3FIb7F+5v+6uJtGaDiAp271t5t
ubbQ91ljuUfD0c8X3accJmeVn/PWyBl+siqMYmhQn7oLGNtmWTP/lt9da3wMQyfD8U0EQYjcUNnt
y7m8IUW482IpYaSBHMiswkmRZNRZvp3lkEb/UPjvVhF6GdH0eiypViQuET0ZkIMWA+T5vDV95hjE
Xe1qWz0CgfJh9FdKYpNYdA4QU3CTTcOewOPmJwlhoywalyiBMq3eUbkvL5bzZ99cCWBZUaPUZNMf
JO6Q2cemuDTvq/rzHXxy6zr1Z3Vw8JEoyCi4ftJMg7MXCe6M4cFBwVbXhSQPY2VxfNDKRnrNtZRb
WJsAPt87mJMawU/Z65aPbEEAX3ep1HkG+Nk5lh7gCXezbLAv1XDiBxDv8TKhc5J1ErDgsbKCfuMI
dSQxHfmCXFwHmE6wyEI7MEFD+DvGCkJqk1as0huYnaKasMoSYiSVWdoyAHTI+zb14jJvk+SpyqHN
OiyULnJujZyM/I/30kcG5ZrCN7sPuXU88pM9Py6eZHG9qqgcybG96+T/DtXXc3yEEJfJslSLkYSK
VLkjNgU8YVFAgMPg1ygHuvG+PFj3ROuo5RnFUaA7Z4/KAbW/BIKNzFSqe65xSLZld7Jx+8h1AtY1
tT0KpKVs126SdTzLjOxAkOmJG7BZN/ukmCONTzU1YRXPRvXzlNqWwkRmmv4HQagVjD6OmM2zMqi+
gpxCoealCl8ELCgem1fY1rN+YbEWa+Qy/C0BU2vee4f4EN+IRtw4N0BLZtokLlPELERSuxrXdvFQ
19d1M6jsazLMExnWd4Ia7Fk/rwA2ZJHs6PdQKbegymeCmBoDSgOgURl/v1E5BntOuqXlySAA55Fm
xIB7MYFWiROYGJn5V0yH2cM9p3wa6oBoHBrg8yVAFHePTf869nB20Ai+4hDkcDqLZXvQJEpjz8bT
sreb9Uob1n2i6R0YHQ7jYPf5ykzzFoZB5oJz/X/nnFfTzBxO6xneYaCezXeVbdR5k2FKXgpLpQ87
9Xk3uX7ij6JOkbK3OqqmXbE1+VDO1Q9SNVDwFlrIwznxEGyPQ6Q9+lBRNM8ttla4aJ1GNHKqfP47
RbP2u73xaW3MZWzDj05VRHJJ0CMqRzZaqPJIkfOORwUdv1qtzphSIP5rQHSTOBjhRrLu6c5AIUKO
Yp6b7mYCxDGTRZg9I2Ee4FImdhhUOSFvTGTg/acmGmob2jiQj29GHYF4FCiPU4Pm28HEi6g0xjFt
1qZuN6kY83p9PvFjhy6efe6spf98HFK5DxifZdLEvbF5Yg7mUIdh+NutvMZ/lQ3+72fbnHmGksVu
XDgvFj8//wcWYyB7J0nZW958PdePy3MF8e9OI373+1U5Ioayot0VAjHgI66uVYyT7AkXoJvaUouG
VR1zleu99STeIbXNCzxjOG2DXzXR49n9yy+TL+Y0L3GKMpO9zzFNGfkDsZySReVwoB4mrhduS1y4
QpGv0NznpqNZS7H9peuJZVWQI7/a8t7QaDt6mkdNjwPLhqsHHTIfs9aze7QXVhXtLke7LGVtSwV6
I1O35crD3pkMsGehnsO6rgPxrrxxh68woGiinZUc8SMofMSCRo5zaXmymgXwo30QTgClDIXaT0Yz
zcXMtku4zFokox7YWwvjWcj7IrjNgo2dRYr3Djn0+86PN0eM11vK16lv0PR6UWBh1fffqdS5iSyS
HQ8Gbea6iHHm1OLlZlPW3D+ce+7zuVj2RFvRbwanLv9zdG/uY4nbnShxk764AzgX9Z00cVSWuhar
kotGQ8d4M8NBF4uGYyR8VIISqw6kVlwEAuJeWgB6vUUmFBnapyvquPRWanw8VjzsgmqN+3+udU8S
ThDTlVZKnUn1kITqKAsRm50ZGUU8YFaMN1ZxGt70iww8y7G9E2d05ShTvAdzj6jNJ+FtJZV/a3r7
VtqoohxgROjVL7hsxiNpIsCuQ03hVZrFX8UeRc4Zz6NZS/gcarC48PWe+OrX2VhE9NivfNcNZ+uS
y+qLlCX6WO/B9v2svNQ+AX4gVzyfoDyle+464IgISeHDyXxIDAlIII5nK13e5OelWPomXbKVxIcE
wUF6cc+SzjY9XyriXOdweXAx1cNp+NtAX/GmQNR3pEBpNnWxDyprKIc8PCKVvEJAvfI5p/wlwODZ
iXLdCw/avVS9/AqVK0IWLZqcvmKUVswpc4c2/Civ6SF/BWPxr5Fli4t1ZBam9bIOtfbAPjNeUYA3
bNvNtN58dTJ/gixwjxkzEwPoDgjOjBQez0nboavwDwXMWjgObLnk09QLRpcnBoT3etLgOmg4mW7A
TsPvuZJiyXXW/vIjMeZsNik0ZYz5p/Y2eGDilu6drt3TSojWAoIH9R/3ddi2lSaT7fg7wNne3/wE
VRCKCXsUJVkFEfQDqcNxjroZI3O8TskyFLCRBRGm8fB2A0lPLdp6vBWMdaWegBlTYZo9F9tOt5Ao
jwQ5BLtdNP9kvRPegH4JTYd9GBRQrYd/cC0+Ol1tnLjY/BM45CzF8RJ/FXJw8Tmj89Lagabp4fIX
oXLFBTGNPqpJ2sw/9LgIq0NraxbuiKnxKr/ICqLnPSNwiDmHYRYfMwunY19SeIPxTet+2LYELnsH
cmW47jRb+Wj4VgRJAJ1mfCIaAf9LpTVY7lfjKO1IH2VKLlHclMIQUdfto4L1/lB1AM2Qu+jjtWa2
Qamg0EJOcyKBvLHNSgUOh7fd53D4CMrJqdfBXyakCFDk5tjpiV3BTMyooxexzm60FM7ctSr8MTwa
MF/7fSJQL0pOwaPasH0+83vPtn9Z+aFkklffdlX+OuUApwSEnLVCeryPnu+4ik8ojy/ER5v1Y9Gs
lK/jiSJICubRPyREdmW1aQ3buKpidn9uIMs+//DQ/K95uqJrfGMh3slDyDVsUb15raKFOdETL/EV
7MYae5cU5G2NvggzujcdvfCi3rPA3pnLkeuxUrhlxDEMjY3oYJhu/eaRoNCKlw0/uu8bzYSXCHab
KfK7mjAJK8Z9ZE9c+bEkju6U5XqKbIi/muXETl9mBP/Ni9NUkmjYv6SNV9DJnMUITO3k0QWJIBiY
gBQB64Bnx79Al8ACzI+pNb1xAm75ARaybVVOn3dViG3IFPmQ6BXDg+Ht4+rrjUOX//14tA0S4EMu
OGbRf/gfwdPD4hZsP/0qlnHaRrylMp5AODPskxUDT55NMAeJRZZLKtSFgJK9xsRmYUDAoX9YSZ61
vgWdu7pyb3bd/YUFPfsrmF+2ephKMVSY1lYRDFbSOCnBVXbpY8NRNJC3yBKi2i2EKrcdoOyFI3Kt
BfhFFuZLJTamS0fn0QR1Hj6CBmIjDXCjK4AyAZUjtBKE7/vKI/b+3zLafrbd1ER2kYecexRXQMQy
FvcEgekPMZ/TMIOZsKSIw64zearuFaXwDDhoPzkFSxu5423MoYrXWLVfzJuw7F3reY9fpv0V9+3Z
Rm95pelFsabtQIhHJqvdOUh6UbldCGj86xlBnBrGAKJCBAEuFtdZVc6Z5o6Qm0ZzjhAqaybZu+m1
9aA43jVoo1yTB5Cb3lWilrfUk4R8XFqlIJdv4B5uT9QcRZrKNfdURhwiZ/p/CVwYyxzBD7fr8Ont
Fjkp786PUvuHHMqpv4kHRMgJN3h+OoJ2LdV114IcxgRyLfkx/2VckTDn7G8cmRY5fcUmuwnOxXxJ
pztOE+Dkwd41O/QYae3iywQ5ZYoTFm5M18GZZZVxJTZ83G8Z9nJvngfSEkjl5TzPe+egMyXIOwHJ
rsY13BaJJ9Ks3ULskLlpsVSUsGmnX8XXmxZ/1bFej4qlKkcB4TFOiYJOHoYpvQUz14pcDZF8gZ1z
cHib7jZH+ujza6UbOBgp2F7K/ot/8D+fWSEqkf32rmLWSx8k8+CKpyZxSrgpjPBJ/ZS6/SwBQit5
XEsB5G8OqT4FFd+p6tJfEkeiUvduNV+2cIIrvUqKxieQMY6IvHv8txGDwTYcbrYZK7J1Jqy/peCJ
SDiAzfc2w8BUdtuCIiZTF3m/+blCZnalAvTZbTpMgghMgy3pDtewj+EOq6HVRZWyhF4cW8ynl2le
j7MLXxMNfWl3f48xVhL3v0bcEdE8kQ7Bit64pm4VQ7wEg7KRZAhXR/PBLe096MS6FBR3XCpVKYDF
DI8XQ9haK2ogn+8KGWl6Tx2yI/2hsa0qJuP9K+dhsLKuLZHH9x+YNYAv4crIbg5LARbBCCMrcWmD
HEN8DTRuDn2yBEUtVzZR/MzmkshrMNxWaLLBPDTNWol9cuFZf/9NjV8qmu+EwJAwZYkaXrqV5cnA
lEkrt8YUgeYWDj/mBbZZdFNbgapvmuDk/ONjKkTn1kdPb0lZeVIWX51HouhbYVj7egcgHsDqZfEL
lxMYm1eD2g1gsPGA5x8JppQiiPlx49tqO5s3RQcyJ+j9tDYdb6pi2rlGT8MOSTNXBqmTwMV8ouwr
CPRdKtf9g090C72gMIRjd9e6D0xKACjEYveYiFY4EzKIURtNyLvRFHXosZQhwS961lxX+8o3S9HC
+2lh7g2os6BaHd2vTJ093DqymL9bnqrzCyl6zqJkx2AkrMx70aA7ddgfcalM82sDAYaa19YRUDx0
HtCIavxWGtxH7xS6qB8wf6sb3iuH7jovaQWO7OHk7kB+s2VtWVMWXtSWB8Zo5/VO3XA+XlcpeVuH
ZCarcWTnJdRtpdzoqDVXMIR7vvuJH5DalmARwJt+dxvLDYyEbaBzYOqJckUHGV5n1fzP1BmDyygY
muqBR+9KnUc6g3nPI6/Uf6j5UKY0pUp3dHpimWfLxJGmK58kVwBXuFjzz6RqtdMw1yuT0w/pH2QV
B2KSPGO7x1yMJ/al8VMo/Brra8+h+AfaHefJx6dZ2KHIbCwHIQc7rk8Kp6IO8k4weWLV9VPisMVM
Mdl4FY3Jezv7fqNPTm2g8RQ4VkSAEMzGYgjJci05p1ap+DEzeSWrXWO5Sy3iuPz3xQhpwBRF7FMw
yTkJCwHO7vrboU+0L33nweHVgJstg8+ZguAtCgpAD4hXjJmVOWKZIojV1XI45buQJFDTXVVSo0GA
MO/YrL+FfpvCI9+O1M4xvn478zlG6ZcBTenx6foMxw5ody1ese5RjSBP1KwQkTkM84tOIZBVhSkR
gBwPU6MsuVsLRL0m1QY6uvFzzsqCEvKIE2CDYMe/qO0/IpjjDOVL44dHtjfSTTOEkqmKQ/uGYDe3
kTJm/ugkNkTMrZu/sKUUhsKUKDvy+rt0Jy2wDTaiRhsTgi6Qof0zPUT2If7/uRPKgJngQx+QBirO
GIcShLo8LIk2+khTt7NMXGMON5Bvx3lca3ZNEcnQCY19v9sgTXwbWfxLzH37lTZ3TxTJvEXd/r/t
WNsj1+43y/QaQhSRcmYycpUbqlL2cRgWALIYxl53C9aGG+5zwtt63gzVr/qEVfFPqtqsFz2NjNGi
UR9GAnqdqoXTWlbXcr9ghDMRu4eEDpn94eQ7Heoj2QY7bBki/CvDckDnoJz08gMo9ojVgQqLt8NI
7Bd7vNf1asJW5S8jlZ662ocvHz8Q2/Yf5+unkmIYVvb8ocn+pwrT0Cb1+v8bOwzj61rrhUNHGiPk
cdnDj6xMV5bPHcYis91PnDyUCUqDGtBy0YgKFz4uD3Or51VnKebTO8FO/T/g8xspcga8j3tb71BG
+Au+cTlxbFR8WvNnEFOwRlhvYK8qpVgbtjfP03APrfeGxqLUQLfKdWsKVkhXf/Veo8FJe1GgLt5q
pDzwVVAzsNF1GfOWY88nvAOQ9o2z0Nw3mzA2T/LZsR+Dtor8iRPef/Xx214zVYfX46bDH0xDM8U9
fPHEnwwXyl1V2hyYVm0HkgumatIWPgcyNbbugf+pD3Zt88u7TV9Zd1Um1zAjsKGSvuoMoqI1S0hC
AzDFJHv5SnfUucQ9bAjnY1LO6bQzhQFaCXmT2QhF30oNhNM0ncwC5lTy2uW1SFaf8wZ1K66rO1TI
Yrv+ZrTrgc438AwQgsHbJ4lJk6pN0Z4EH+Lu6PKCeDfbYANGaR2te3njXMMOXdgzly4vBc6TqYEB
EQqKZVyah95C1uu7viEvp+YNDnQsjsIoEWVbNuA8feXz6dzigk0b19icCpTOkXbI7Z7LK4s2o1B/
0ci8bTT8oEglXIpHcQBQDWM5C9LIcQb4fAtXc6fv/6rOSzwZ7mjObxJSRusw9lzji7P4eZQN7yLf
WGwXTZKKGZHXAeZfj359hgyn1lgyg8zZ+eXL7zwUK3YVl86vvQGvyOS8VCjeUnZEaRI1VIe9g0yx
1dPTLLGA06si6+HG9IRx31f7OBWVITCrfHj9CIRxo5mD+/tKFVmYl5tyeXXZWjyPyttvc90PF7yl
uuXFQVUTai27w0emUa99IJU9UPifnw7KFk1oLDMLJ6w/PCbxWyMoFIghpf5xwB5urryOLYnqbpY8
ozBxbmP11Yn5VBYryYiZAFEz/AZrgge807p3Ld5lRYlI575ky4QXpE4abmeywXlfpK11HC8cAGza
hVRWRi15A7GNq2yPUzx2wztcmLhwWqb9LG07ilUr04C++CeQIfau94FZC2W4xU2z5BmtQvRcObn7
z1l6UDPqOrj2FaQ3SGUZ0a2Fom+rZiCz/RSbLLC5XhBIoTr/qJUy2vgryK4hOuPcFCHwXmfC3zLm
w3VjrAweAZ4Vls5HdlrBejtlDwFgSP6sn5bYCcEPs2ArTTaXcxx0guPA70UAG4SWj+p1xlnj4zbC
qa28087T0517GwYcDtkuoc5QlQbd4pnYye2Dlzc0oBcqqX1gYru+/CkS4JbRHu+L5FoyL1uzPGDu
EyKJRGtTZd9ctOTCRUjrqLyevvNRlBAdKZ6U8Uh21QJC4MiFxkZ5AkG6ErfPCjxrf5aREn0y8abi
kASEj/ocwQMG/zmWLJOJ2o/PB9OcUUMC7T59V7uSemkSXzuaOEtMcuQh8U1Pk70XCDcRQudhKv0I
KG/4VYfCEOa6O21j9KymhZc7+/6kYyDRU/XgrFyNe2yXaG2+luiVfQnfT2A2hCdkKm76jbYSHZxC
Q4SDiEnhdYRZ5cYhz6KRaHItiOJ6+7hPV7PqQrbxPAbWclgW2SgiGbGwaxt9D+J5q4sIgTCUs4wg
R2EGC5YHlv+EipyNFNUN/BYvKoCzFpm0lpYS3lBAqpa6Khw+O0+HS8WNLvgp1msuV6GqCd/cxpQJ
FJ9oOzDiaueHsPPXwJ3snWuo4F7Mfs+SS2+Yn58CQtRNPNyKvWnXR+wAtTO5khNIUrpkkztpJUgD
o4Ag1XTLQYdVbr2fc2NdfjYREfam8IJVaFvr5K5mRZEqbcER3JGMnuFr0N/yCkxUBR/jRTRmFWSA
N8d605gK7A0ecpYcRHP7TXgY7T4eKW6xA/CM5Xh8/BX/zQUalk6KxdeNUxQ1vXSymaNPUE9e5X5d
f3SIHk/ErpbdQL5ojbB6/eDkvRU2Wh3VsAVW53nBoCD3OIcacRGFHgCkpwH9jFoQ2nLUQ6ga+JVJ
VrRPqo2PDvCKwBLpCrMGRayjMb3ZvukJOuPgwCkHcXca3Dh9TvnS8vGYrnHrzdilzK3e/4dqNz5X
YlJ31csjzxYEnLrdQDWDR9NrkCh1iRgkEOeTQ1JnUqABaZd+QZ1gGlqBCF46UNlihgPRI6svsYxr
XShWyqnfPMTysNyj22Uya7+98uBO6TtOrZqD0tteIUw/EUZMGkLwRYVMBg2+OCDiXiuwGoUpUIOc
X4Nioe1d5JIcRBGSvkgSw82PjFvdluDmEJG7Ue093vbnxCI32kCN5yZ379AagOITtZUwplqsL6qZ
sdeiP/JeX6E/kDi7p/eXB4X8/PZYRBFW2hYPjePpcFRhE2CGk6vQXjiFnZHtwtTVZ0cY8Fuvo3cN
PAsfROERZMFpBCE66bJxspy1OGavxvCI8B3jivMi1PS9SBWifoK2t9vHr1sF5ppfsQ/YVFAqlOd1
nIqdExGCFPOGNFs1kXP7u2ZisUfA8ZUhrVTQQJLe8aYcUA0wc4Ntba1c3RfDDwuzTppLuo+Yz1tq
0qMnvjV+Kv5a1t2/A8n2vSVxrMjLJSIu1veUee8c5EHGooGZjW/nmiRSkeRWCtv6cCZKcSWUlOUC
WxK4sOhBEk2QeqOIutk0byfLN7/sdBF0Cwjrc00E0mfQi9lR7pF7ZtnMnJRTaXj/338ljkMZJ3el
q3BCUWIz4331AM01gbcxZQiJJyZ2aKgvKLCWphp2zQIHcj05vBVj8aMGbqCbIVsp+v7CYDVGvivH
A9r9YWn/2x7P3HO1uZ7lAmvDsPUfyPLdEagm7wBJY3GKGpFWLgJlyswm9EE422NdXmNTiviDE0sx
jvwYZCGSE2Q5WphKwAFiDYoA8v8s0cqp/wD8JoL89IQMD0qGtkNlgZ6lskB6lh2zPdrU/luem2A7
RTVonNpPH/Ha0Uhdd9N5WZsVSmFnmmjraGBFm2CLtYxWZ8irnVkgB4FiytxndvKE4jJk+lMP4P6l
HLfbVaOOvIj62VRP9FKgbdRKjhKj0hJWxUf/VBEDdmrsNUp6+esiwSmdJXIsaDwsa0k8uOsKST1v
+2m8/zkUu7wgdxVtH8OfysQrc2nNg8B2bqn6t2gNHdPQtvc9dbh00ms0RdvBW1JPbJXY9lzT1Mbx
yriNBm2TrSrSIwG63O59mu31gSDcB2ob99znkqx+EAgga5gv/um/S7t0qupwstzhMdisytje87ub
DqTfElVsEJdZFmdL/fhI1mAAhnCOk7h0N20T2A2/5FFqXaij4xAIxmRnu1cWROKWP+vzNXnHOwOU
lwgPkyFLFFPeX6XDMI9qYTfUk2zpXJmqvScl/bzh3IUWEGQcW3Owm/l2+YYbXptkCUSG7iu+leBC
wfl7qE1iFg3GJEx6tt/Sf52O+LJERQi8K02WYY1B8+SCGe7DfE1gJ7O+pjLcBg07TYf9ZWqMjKxm
wT32/7pQyAMyZW8s2/ruWubtq/lLnj4azALRVI5np1+rPGYUu3X1aE/n/Sz7ESYXkmUDdD6jUcRI
xPHP0Dt8LDKz2GwRGtWxz48cNxpMPdMmweCsFaFGleOk8lSyRANh9+GlIzLxgSDCG43rGbC5cDeq
Uqj/T1H/iK2E+Y+wxoONoebO/uvUlJ7sJIgyPXAMfr/ihyl5kLNC5lwp1KGjjHPBeWdqKGwaiEux
4qg5CleXzDh2vmwbdWFlPqd1p/1HgQh7ii8MweJKhyjWhw8vml4ncS4bPoBQ1+bmUHXOERobxwMQ
i5NJhTC0gH7yvRdFm1orOm4zjcahQz1rjxQ+4T0D63iKnlWU5Cd7eQ0Nmk/6oDnNPN5tC+XUitWH
mC41wL+TpG/zTR8rEDEeVWUBC/SLoshNfyUCZX91FEk5buOOHz4XrQdUSTT0ltuDuF9mZz/g6hrR
K4SfrhgO8gAaYtryWCOGEdd0gFtgKVyPDjCkXa5Q7IVizC/MATJ9WTWTet4bEvQUtAzDAk2VBJ/c
9Rcks5gY1t81QaLWxyU9JoH8KaeoJdYKayb0OEDiuLYlI/LueWVpbsr+c0dcB08bCDXyeXPC/CGI
bdGhhbuU+5cFSnAR4c5hjb51NVLSJJ9DBoHJ6V1h9/8oBMj8PKig1MVGdqSLNgU3loGE23QFBSHl
UXotBDCwIFhoXbPyoWDfNKYUZByhjtW+9uymNS7Z2iDiM2D0xasNajEfOP/6csHhigDJMqmWTdm7
oLPM5DcHDbplddar5X1u74E5UgsUbs6eoywvKudNDxzDng3f7pXokigb/yJ9EzG0luuri/N1Spxg
HRMNq/nIsoVq7Niaa9JmGxejBR/NtzGNUX/wad04qFJWCwEW7uTWUGr786iMqpyZnMORlhUA9UID
Rhxn6CZfE7uOa9Yo5E3P8l7vSYu50VEJLE4rgIYoostdBuUiAeraY7jsu1Sy5oxUaLJTYCPTtE7p
ZGkrf9K+GBkhcBYSy2D1FCmoQEPQ0oJaNlhsKOdmc3IZ50W5gicZz0RNsotKAzlx+DCXsWe2dN9j
lGZj9WLBJoDFZNmXpqDbt6O9KnKMDZblVLsatYsOIENwQojHRfk/6Elo5ZdaYGJt6rOvW9wFLY92
E46s2/wIisVQx3CJL32oN0eLXxpjICw5j97lBJZP2LR9VD3XWRXrWz8a3dXnWs4iTaqfYl4t3uC4
SotNicppm/uMbiOYV5sRAb/ZOHMU2EFjIKvWSL9VYY7zN+FXJ5tkWdhDOi0O8nfcELdL/aY6LHlr
tYd6csKnKPcGsN/jEUWHIE0+ET7U0+6AZ+GDzuwHycvWM9xJguloDdi/N2CRkxo4U3UaNMEIDo79
EdyCrSkvEoJCj4DGYHgxj8WtLuDDHT5AYnePS40B3rNC4rDRVGqeMuMpVrc+T9jkQ6j5EYowgvbp
FqjPzqTU75JZjQRuBdc9ftzSfsLB2LQU+KjfGFA035omTXOk02dd1xVqhK8YBzrwrTINbS3Wo77p
3tKzNt0HLT05AykUtrBT40GkjZpZPYGcqHHQSWqG8JvnvGpzNLVelSpo+qVYCYxr+8DV1esYiV3f
nYgY0Gp2u3QkVV4B6H6psWX3ukYDZ9qNb8klmfzWWGP1OdMB5Z5xd6FzsuaxK9Dl4c5XGgOc4NB1
qFI9zwABLyZBtHbdzH1qFuH36juyzTVk7C+j3HXi7YsfHZl/tOsNZIkyXxykgmx+uLLm2Q7Y08Gu
49MzMDAuDrFJ0BaSFBXGNw0/mKIeuRTJ94VIgzB7kD8tDdsgP/7WPzd492/3RN4xYaPbM4fdeJB8
yWSktyCRv4mfJH+OtcNQMQDt06hA/AgAxoUuGu2cV+qLeTjHsYfzXz07Lpj8OJuh2PQWgW54MPay
0+uLCIbK/mQxDruq53SMrlrid9huqAYe2Vi+DjDTA3iwJAcBz2HiI1YfCxT/TDdEpXIioG9ydEve
1AmUBl57pYmyYHpbSHfQtNdMsIN/NPp9WU38MMpBX/2+/Etn1iOdVgf/hhIMO2kECccRINRPmFbN
dzvX4nBSYsGx4FuOO4uq0GTDqh/Xq6snl8kwyQdnR2ftQWRGCry73wmyTTR4d7kffrzDjkimhply
4YY1hFh3A4zkz2yD/A/keSOGwfY2NcA5UYLzpcSMa5EaiFqrriBtllqb+eyjur+5xrWGkZ2Lk/aB
vhTpQxlGexYnLOP9Mi51N1yqWBb8/PHmAlle+M4seXX2gCIE2l49kVJdpZXthsBvxrtmKg1AeV6r
5ghLFmVQZdRZ9BW+MkBgvSAMHzy5hUDEkhGskrZ/O3TFUlEz3h+PStq2u57pNr4WANw6hNVr5sLm
m0izPYxi1ljowXov+KzjPwSPzSBF4eERb54avnhSb3ae/51c8hNTfx+J2rO1ZZ9Y1RxAlq2p0373
1BV1oo2EcLg78UOeNwFLK8r1t/ebWk6aC9SUFBSfJxk71CG7RTbjMUwFAsXkNLI2GqPOSQSwfGA7
faU9vRlMo38zmEjlBjtN4RzLEH2X04CFd0GujW69VW8GTWwDQJiElKH/+twfnZpY2/I9523S0Qco
MSbxFg3GTLYq2tZBt4pGzShQOyqhtXLSfEOQ6EQ4318QCms1zPlfLVrAnYGSXK2bLo+OV0FhiRtK
P2CAU/7zrPKoZF097yhiMDD/n+EM7gin/YUExnS2WysNiBzsuFC8Mg7drRnz18/EJrqZX6G5d6qX
McB2GDEhd811Z5rQ99UMQklFRVyQgnyuMOaO0/iuIY1BXq4WASh4n2nK2QiIZ38BgaUKVsC7cBCH
axVXssi1BcgXEJ9lffMlu8o+EgsZbtOwcBlVB2AVafZPD8ZyFYGxCC4qbM5W+9mRIKrYPGTe7BN+
3zp8znGyu79QYWJCk5p3PbVAxrecsY+sRk+V90CkY8w7o7JKBV/YHZhoYiukEIFQEr+LDptm6TTA
i0TiP0NzO7bSOZwByH4/NpNCsK0qO3sR8LHl+t+KXyDzx8vpm0rPorqtDsnFV7P71l0WS1+Y2ENW
N7LayvtCMMd9msDo2d2e31n6xxxz9BANNSo1sCTEJKx8DoxXQzAadRQhE3RETjQgnZVkvqAxJUxv
DVEMsfZrqEVijtoWMcypvsF/cI65n0jUjSVGwpadhqwet+daoGsBYfxd1erXTmIaMP71x5IF9kvS
C5i5riRlqpjMYGy5u+0X1P/ngnvW4ScuBocvZ8wSVt/NYNeHg7tEgh7eaI7LzynojeB5iN5DN7uz
lmY7M3t5T7UA9c1k0ACEgyCsbCxGddPeoGcUvuRXRwh0UE639zr68Pfrvyrv7ojpeMG7FyyKaS/0
6p9sHIgwdc7h7oRDsm3KeVR1nrjOd8gwBN7L773tvnTOZLWaurqfa92dpbbTLDXzu6vTXz8io+IK
LEawB5VhvI0zynbr5fPzPTSdva8c6181idQU3Ih5DOrI9vm2CJSVrDRX8fXc7+bzzq9A3EJRjWZN
7L/JTTXMvsqfwxZKVzn8yJCHr3SWW8LWiSp14INAcR4zx3V56VHKx2TBZsz3W5k+UWceY2s+Lbmj
kDfQojKFIBZKYbFL5GRyoPe90CZf3v03+zgY7netnlEPkeB7zMg1aobYpsnU2TbXcIjwn7IJjfdj
Wvx/0LUT/pT8k7Iiw9X78foxYC/iIvU0tNOXw1OLFQP1D6Y5n2tDXGeDr/CyRVJl7KeKNBzmdQcm
N5vRLANlDS34tbL2LYeHyTU0iU3JS67r2Drsp+NSHeOn3XfFP3BYSp4Em0Vg2RjpAv98o/5SmM+4
LBH9JbYZZ71awA2WD0uDGvI0GXec9Lq7FFnrJz/8Rt54T0/1LMRCPPZzVveJwvoYuo+pWqhqwGBd
2Y1Hk5H0SuHX7ELi1VRcGy5LGa9kB6X4ap/kYh4BN5o++ClkKAEWJNb3IXZo+k0EhIbGU4MIJZch
rWV0ailNRTB92SLiqJUDbSaAn+prsyKDcdwz/wKku0T3f/YA71Owd7w/aamNoVBmTNKZljoTafk9
H3KPdAyqhgryg4uqiFDHA0bbayGBvD5j0mFjrfQXwNrq3YUAb2axUqQA7Y9mG2M9kKHbnuuSX5rA
gM8E+Sbb8AmvwbwecBJMLeLA0IVvRqHqRvWh/eU+EwaM8c+GK7wOsyTdsdClRXGyA/kXbTegCPoC
C2QdHf7HdMCXVwb2Xa56rcclaWYGDnb41elRXHnVzSimYV3VhPuoJUumH9IJUiYj5hjWbIwQPR55
pkWngOiJdgNII4GZoiuJ0yZVx3LMRveXdohu7LdyosTPT/Xdg2JpxdLZUiN1i9k8vZ3+d3VRNGu6
XFkgmt94a/ulYrUdURMcHgVmfvM214Aij7WqWmjJBJxUU7p+BWh+iaeEwVbMLCeyv867KiZgqlF9
itVfEg54s2nyy6r/HoY28yQr8fn7g2WMLxZfm162wJLg1uww8kSNPlTOJ0p+uvAsGwZZFstY4cGG
9m/HA/bfcdNBveOx0Y+Poey+nXoaztwX9/YbKtfx+RUr4gwj7rIX/EAghXBMVxFmNqSNwYMnPwKA
8Bq6zx4phxXLF3aDoyElFr04A4b8kBiDhMBE/JkOxLhl2fPzLu4Tz1EhfTWUiWRGgwpw+NB6xTky
aArn6Miu6AzdrYmOUF9KvQ67Fap28niGz6OCSxC25WC7t9v/kzrFh/XpT8VMaJ5tvCtxnp7dfTOU
FjN5g1Zc3d/Tc6NtxUO23QkA9gHjBcAywyw53u9FIzMMOCVpVXdklJ9CQUm6M/gVsNN0fo1Wxm4O
fEB2hyJ+cyhbsfdWBrU4q0ZFm31xPfUTyH8OwcyxXVIMDGiMOceyuHxmCu0oqDKTQCdwYJXqtHSh
uuUxel45E0hW4s2Uyv04WWdsGlXmnXIAUap5Px/rpwlLxCu446anhK10SzSfIcZ7enVgqUjyLybm
BoReMPBrkX0tYewEj/Q3NuM0y/4dmuhStx+t644818Hack6/rH/XqvBZ38KtKNbhuf5QUdGg3jES
n35jZoB0wnKD6cG8YTJJkq23FL5FPWdh+vM28XMKRqRnDGuhT0vEy7TB0y92T/SmEXgAgL4pwHWx
Erl99CS0ozwHx1PBJk+A1RMMygPP9jgus3JL6wIasPufsmb1BSWgX8aqoMk4LSKwljPnhBZYd3vu
2ndCPMp3GRsz+cQgmNsyXe9aDOs6jh/mvXmr9r+qiAvI4qhZAIsPZ5zZ9QfepyL9dC7sQt5nZKiC
P1xm7QKG17ZJVt1TxFC5sVi0kniWV58awzQAy1QYoWXWP2Xpd3Hy1rzqsvkBXL/gO11yHUgPwIS2
QGg1/YPvwjzDHXndC7bodd1MpLGHnvksl2BNE4yu+nWMJ3bIqalBMuQVrHIMNqBUretQ71lkJmHh
QpjzDRYu5VaXISEKTPloapcKY4eSk2kLUyGIDCqtGF68zdDapFHubcKuGCg5V7+0a6qtZ/STQUTY
Czy23ICftxaQfUtCbxFduwc9YAJFobc1kUZ3zDiT65RO47M9Pqb0f1AHoX8GEEOm094/T0IGD9hW
BbEGvTqh5dokcj3hFb850iaBkPdgEvz9XYm6+CEFbWOEkQVsxbU2RxiJkv1NfRXqhQ0wkUNrHsJ3
u+ZjkreFNwQClnGJFZoDum3jH4loklDXNP+mUy3xJw+2ekLd0xt9692nfC7EPhWsXo7bTxHMkvO/
HOECDwEPDlToWDaYXzyL6RHgAImdPJHXbh74k414CmKraScJFQIVfhQEbhKN0bYk97RDLvcG+oaN
0sclkogO6wGYME27gaGcz5u62pjn70pT1Mme506CSzynZKFXr11NGyvLtcVTpZ3QT1x3/En6ZuhK
aEVQZ8EkVRjBinMGRgasPvaNJWvkurBHvI+ngkHLcMtJ5Mupg/+zHFH0ld2ZkT4FSci8ll9UNwQ5
1pflXPG7s7SwPT6HCpgmfeiM+1GZSV4eSjmnd1v2UNs/xwe9LSLkpCGY+lBliLXs/4/P5rCQA6oB
LfgCJJw77anOQ0708XaR/xAKmG4AyEOeEtNn4nfu3VjV2RO/0+qt5Kx2/bsL93VF4gVHA8pxRE+i
O9mZDOIfYJxcADzQ+MUsUuHz+0+FAbQY23gyb1xN0CKrP/4XVgozvck7/9gGQWBGUQzueoHpsNKk
ptdXTHitXYw/JvwicBjPz8rbe/GwdvzmrGx8KwK6n1+FWB6pA+25h++Uxcb3IzhFa5CQTyIs4NEb
+Ehg4pV+kd5UKkdwIql4p8ZVSpcz73kirCmeX3Oxz66QAF50LPHfjAgiby1VPZYp4ZIjSLwac12U
GFZPz6oRMTzjViaSASZ838kDxF30ZyCSPrX2i3k8ylsoRbnV1ug/0hbm1n8Fb5hlUCtaL6y8z+Hg
34Mef57/2wl3ZUq7qUHmZXpbrOEe7m078XEwyOPixAh50ioFVSUwVU6mYYTOdEb6W4KTJSnhPYPV
6bol3woRzWoUPymf9luN89REk9CJcG38tnBBtk9aiyLXPHy7uN4qhuPxN37pnzuW9gkfZFlKtIEK
1vh2463Qo96adJOFAZmTpcNq2gccXVpO7xnmvdAmQvqGK89/N+m0e/OEvBmBV5FLK/t4k1v2zBWS
35tuW7flu3BnVDeBsbOo7YVoj/pA/h1vFDqUSmt+9A5b/vwtF4oDAKxgt65y4NQHPEQp+zrfQStI
AmFmlLtrXDKQie0abrW6WVYrPasT+V69xYPNmz/NJncvq6wGItmwke0uH+nGdhzlqfAPQRHnUmIl
8hx4IL8gWf3fN4G3Dx4VdIbpCWxE6RChsYt+Fe8OM9q9GL7urFuMCF03QyAQUAdYCGVPbL9nW0Zb
ht9XS3tcykvSRqZnymXZbuFl/hEWqsPSt8ucBTxeE/D1Iw1qNc/kWOKkgUVAHuf+h2mPkMvgyPvS
DCdD/E9A7+cJuGJc3yieQUcxa25+5th5fkDktrDnEUfRYLxeIhNoeLVsjjQ6/e41Kk7rDhENJ7rj
mLvLFTiKSxFdJmb9QznAHMGDMp7ft3/dlxYb6okQBnhUQpP1qIoOW2b2G0yn0H42UHhDi5ymkEVs
1X70N7HrjaLnunNhMENBl+kgabH+N2bm+8crklyScPuDSO0vXOi4DjnhXJHcJd3Z84RBSOmfu0Ri
/rD/wsqUGG1pLvKEasJ3RAU2HKdusyTeA+Qqkk1WhGcVqWJuxFenW6hK4Uf+kWbU7SGEaABhEb+B
k+oU8qsnnPcn0fcanOQFH1X23OfAjXm5qg5vuK3MElXp2L9SLM3vdEL17M+hlRMOxsye3J1yppLr
YeUnYYdkM3pUQSibDAJpZcsjnjwgjcR424W3Qt5C7JzxzLoj41sYG9Q9eGfH5BzkuhQGttAHsJB9
FOQmlZJ6k+QB7LAwLn8ORuxkGaBYpd5dBjgj2nGmQQrfJrxrT4DFiZPPL37UiZ7mcjSJ1tqJQlJf
Ap5ForVe9iZCkew028JyiFryrQdCEeD4o09OEV/NsjzbjHRMkzN4BMjPZRplI2s9e9D2Jco8Rpm2
3EKvVWc0JigpkiK08AjO9PJQMza2D8wG88Z5wL1CnSDlnaJh2BBwGt0BuOWYzADZ5QWss3TQfWmS
TAARMBtUr9ruTypbQTrOQVWOv9ica/yFgQ5EENPNm/HYY6w88JjM8ScpNLuRwlgwKX0HFyB6NlBV
Py16AtVWJaYeMUosJtk9DqwxImwk83oSousEm9nf+k+fjqLAAcc9NWZn8lhm6s8Z3pXdacR36Yw1
edHXDe8hohUOeabMcztSvfj+/WOrbwxC15Zq7WEcdQxRzfpC4heC1Tjy1z5TUA3Ji5lHhybrnAOy
569H+QYunr/wqn9v5CwjqyOp4TcQoc6gF4uK/EoIFoV7kBcNpq/5dPmVVc2lKaiYX7wdTqDDAvQg
0YFQPT2n2dzEawXam2iQ8QyLPRZHLqB3TsO0ARvTQpv/kEEYe0rJ7DEH32l0F5j2ymjVp74XWW2I
pvv0Nwd50SUxZsU+2eC1ZlDjw+gOb/D/stk6BIoNyKrWlzq0lbjNygt5hghDUbBhrkswYgxK+zOh
T1PEfpY+d+UMvaeXRUqUToJYy3hDVKk5WfTtVa3osfji9aWEmbGjmdDIGvc9S9R4T7oLx9aesUlc
SGjdr6S6Udj9mOX+d5BFYcARZOwus7khDM/kEkFsd8/XmcmyUe4jhGn755Q5ppfE12okfykkGvt2
U5BsZ09ubTJjmORwjIDcpmlVCjBzN7Cl/H218HkeFfIesRwN3nWIEkn4yISdEXzJCTSVymqH+mWE
LKiVGwhtuhPH5wackBxPiN3qDNRvj6fNULLCEISRb5B/Ju7kLIA5yyAY4F4j+HnbLK0/wlPuEJrZ
19U6P75N1M0oVWHOquvAJaSuhICVsfIE4jW+2VtuRKDgloSM08kHk58ncXiRT7MBdwXWO4OPr1q0
BSyO2E+1ov7Iiy31eDfsC96WbapMsW3qKuE34V53lU/YHLCthEB1NC2CEP13v6N6v4URHmM2IJCo
9QWfAgm99hNnfUQDbJXzrLJu6z/mPt+f7lzurhRKX3rhlUmHsCJPIhZUGSAExueSQuCkrsnEokyk
fCA5XfW4Z0GeNndjEJQ4k/ZKD7ZcMsUHLBx3shSod5B7LWMdTSFQDNymAkE7THaTkxhv8smHWFDh
VJ0ZAZtmwUwT8EelsX6OJFgAPdGPD9i/mAeV+0kB4X9Vn12JQaF4GsZKYHZVCtSc213yFnJ8wUtT
mNzwe1jJF8hHuvnYZT/Iul5myfSR2/H/C9ZjfLdl4muKyKvSqsGaCcedzFxOk9Nr7H6b+/9i6l+Z
su5DJ3V+Z3z5tJbgZ0jh5KNZBYnHCeGCkskeRzRWu7fbH7+IBTqcnsgCb8G6CNd/xZ4jbIKPuVft
OH30G06Cxiv87ykOw/dfY04s8q0BeX4130d0cKxNH8kPLaMzBFvgu/ML2VqCGPNxly7fEOA/ue2F
MlS4T0sjXutlJh7puYmZvl4bx3q/UZoRVJ7AB2wiCe/OamG+Jf8SK0bKs0LJSUCKBB00sD6vSPxM
VqP/MfC4FdVpz7jIOoKMkWxv8pkyu+H+cSQkRD2RwT7FFpkP9QzDCLin0l3aLbMDTJovKjv4rcBf
EA90MsxK+TtSbR2iyG2CxQrpEBdo4Uou0olrXI7IzwWco7+OmBS+Muv9T1pdvlLA+nc0Ym35fBlD
9ABrH1SYKGDcOiOWENDCkGTkri//TqLYIEAPRq3q8tHRFS2i8/olRTZG+0/NXyLQWwbz1wEUZppy
2fsis8U1cvsYY+WhhuNeWk3Br1OP1PklR1G++02rF7gkZ4YhQyESblp8UjesD0b58vtPzBnWeN/H
oM2RpOTp4YsAcjLhhwV2EabfiAkBVSXjcciVNJU+iwwIxZs8kWaN0SOln8dgWNi/V7PBOPU8oFPb
PbkSZQvm94fjCM7LitC6KYkZLsvGRYb3LcjKSEH6zQ/hBRJnHEyugctk0hKAuoPP2qLLWMKjBtxD
21j2Fq8DgDW2TvHzJHJAtx1bzcHTOhQukSf+CyDW8WxwlnZj3PhAQ1/E793OYHwc2lFeG9pNNkzF
W3C48k1o0rbnuVFOcWe9q3UzJDHBKvXDdXxie6d6RZGnBVVczffxUKIjXQ/NWWPAzM8uP5lV6NGF
BgogHVA666jLGWoEKa9dSZswyPOL39aGat3wk21F8GXxFoo2JQe4O/eHNY4lQk86FwjrVrmnS87T
DPCZEgca5o2lHJz2edVv+sltzBsBBsbLx+6B1+isWi5T1orJXSy+U+wPX1O9eZMKangO/gcu7HjU
N/xPmzXTlwco4FUupUmJXczc6W4rOXKaIcVUj1N30UZjpu8QsdRJAjs+EfvKkq+Rn9iVkBB69Qrb
sTT7+X/kLTFNcCwUEj8cAxZyWcFNjYN9x7+t/MWCbMReJoKW0Rhh/pN6Qe4GGYUlceRHOyx5h17f
LHqjGSUvw7Li3TY1Gh9N08HZZbeHYfNaaNOxIJvNKjNUm75PtcOi2KfL4cuSgARYpp/dqXrPLuM/
/pZUVxwUBVmx3jiYtTJsLsLA5SyqyX1Hk+FFy/eFwIxzoJJfvgXGie7OtJrDlDoI669F6QBH6IzS
yMTJkFJdipsjTcdKZfaWVsWwphIY9ofIpqJ8bWupxYkyJWbsi6IfLgJMDl+DXCxJdKIK8EqbCp3q
CVlx6gn7ZClT28sVq5Ni6KwD9mS3IbL9hizdHrT/9soCHX1bgfPWh8cr7rPTzbQ+9LyFe3t3QBPn
705IJjas/GM57O2v/hv40W6OKdWqIspt/OdmLJuDJoEcfh4nmqT6xK9Ii8HtXaErEk2QB5s8SnJm
vq+uqBaR9BXIPWExGc9Pq1C2ZR2XkTpJriMAIpbEtiSbVhgNXyMWg9Uji86kxjOMqktHlBvTzHa+
wpQBDZWuQqXwS0JCwAtr+bIRTZ6jd7A/A0zutMqF0y+MLPTSZnD66fsCEAMt3HsUUTtjGOVKFb61
+mjhCLaeIEwAc8nFhNKc3VGpMuaAnW25J8XhuTXTpHGaLKROSa8ukOV9tFRLN2KHXKbI369ySH1X
H4Y1Tqt2INGubWzjpFUgBerrlixs/ko2iww7E2gC7NjTd2QzGE/B+swRUcjLDTq2VkujgLadrlhU
Vyd7T1/W9PPEQsaadsAi2ssjgwnK2TxyN+3L7ObIpeiSOtAJuL6Bs+c/4NlQrNRXFraFF1ADGNpi
V1z7IaknW4GRyNgdE2xTZ0y/RX3E8opzOcIoxz8ScZnBwERGpJTEqebmXm4VtljCoI7M30JRDqFx
XTXGd+LRHK8963lUhxgHbCy2uRVmDML9VofGL970Nox9JMTU/M40ioZFvhaXJskcjxEkb3HgKr7T
Zu4wTtZsRPkqliJB2pnmY2/zhnyS+SGa/6PoVPmDQjwYj+GpuZY6WSCNwG8Rm8VFf03abYO1YmSv
Mmu+DVk83aCcZ01m26AHTp+ZweM8fbCd7NbyV2mss7trn56LsqGFxQrm4WJkHCjrPUn1WXH4TjdR
to8YOUsE1UboA3DeZxGMeGFiHrStxGKPqJ9BYyw8rqIcvq0YNPJRpuvSxVctvUCKqpthgbL15az9
pjPC6h6oI/Tq0lpYQg97U66CMGsgyudoG+dQ0f0TkQJaeOzSAHi/4BUwc+vbtr/42uDejr12bAfs
LB/Ucken21sx7bgz7ZFh+nQls026xk9YtQFM26umMoONBpW0VHicjSfsfaQ0Yxz+OP1sq9FSZph4
0rt3ZglXpBTL0bufBKaAfDnjK52wz2pfpmdvTsJgjCYy/62hfQSvQOcGtsE/z4pb949C6M/KnMmC
xB8VaJMduwaDEyX2DU0KilzkSNSDFGVlZYorr82SU0Y6UZjiPwJDow/aTp+4hVOeGbx3uDrrifiL
gVl8PT9Fuc8u282vLQKlDzYdsvL4FB0ZVI4BzNMeJsZfKchhZ82ZAwhN1uptgJyP6oow8iz4CqBM
abZlkWUqFg2OFR6n8cZK6LmT4rfUTF9JL/mk9/oKweXfwD7+5vXY/Xzsa/NAr2fBWyNHIOFeTpkC
2+S4Ify12HYyeLhivuf3yenFdQCL4+iIf0k0vLvOosDgPgeX4Mz4V4AV8/IhrtR8C07k4M4qc/XN
IceW0OA6Dcq8vIIQuzvO5o2+DcAlMLve83QF8QY6COAljuOcNGAREtjn1PX8UR+lmfIOEtCqRais
iO8kIv8h5ikcWMiWebX2nN7AcxWJsWKweypCt3TpFCToR7Owz7LjNNTsWFI+se5IKL4DtiBVLjPn
dGXAGSoUxxrVM5SC8T6SiFLp/EWkkrN1F2SafSnaZnA3Pl+xqt8zO8DLEGLgVfakJRnfbHzy3Ofa
kW5OSTmlnmJkBSYr9rA/Ki/eEfaKo70HPMVhGM6yiQTRZM/RgTzW5C0tkgq8FPFNDtJotlnKdbYd
DdueOPHPAL2Lu5vdkaCNf0+ciqxgt6W8GC1ysM7N8EM2s54wGGN/Cs8A2D9bsNKS4XfC+4sDNCpU
f+nl+I7nd1nWtXCHzjyTnrHCF7mIQ72I3FyIOCHBeUkylsYC1QEJl4DB+uziM+uRzmSAQ4PjFbg4
7SrL3KybEq9vbTMmQwZOhMRyvwTtujjJNF9ZJ2k4Bi/vFnnc2Tb+DEkC5EdUOBmpg9+whcy2Ocmw
FBw+IExAlzLJkFzXpQS8tSThPfRdFUCuLGxX45AXLwTzto1xwKYHRqVV/zNET0U7TiCeJ/0ze6n2
MbvTY5w2b/IhDYBoKj1kk/6Xi35Mf5Jbkb8Ri+aoH+X51L4Fgou+qpHTwHiKxt1BbmOxOJcLC6kU
DoGCxzAsx6IflrJ3XkXYlJkdTyVdwsKwUQpcbOBSv19x1o/ReVaZ7KcGL3gYNtzzN6+k0yce4F9+
fgesoelAvORkjHzHvbgZrFtjoE0X23tCspK8erdnua6LfqnvTw9XeCHTvXrb+nvOf7XgILOaCY2n
IX4I/Wbt9poTEXEgwVwkduBZ0cltyj6hrGK2TrPXVdt+l4VQ04bE9z3MvBeRxta3hPbVTr5Oi9es
4wt6tSGqpmX1JAB891Mi9HPOWff/aMRcpCNZo7Nw9Pd5nUTGe/M3CO6cF1yPcviEN+XOLsHD6PMj
DP2m29shiWrJIiUvOYr+7qeYHv/vnr0a+7vmQEB2IzlnSAR4himvj++M4fMAzn15rFN0ls5y0dqN
Nu1nlz9DcKN3rOSaxi7ha0Z3TuBJpKdKE5ouegdb6gU45EwbcRrcwpl56SMz9trs+40Y+gQ9j4/E
VqM92LhBvso/39UhXDE3hxWL0dzZILjbA/e6ISMBOyIIzu8FMWr6qXSyrj77pvK/ybdXOSxyQwf6
TQCUKo+VOdQMJWUj6QmuTxF0OFK1+X3kejLosyz7iLzjnZMk6s0Ynp/BNHY+0mCocpQlASWBRT0n
uX75WTmYbgHOMZBiN0xjQlnapRRXQyU2m4kH8Z9wrhRSJCUOdgwcK1Deb+BhwfTNvwQ6QJBIjpaT
e7QzLKYwpF3gEYw1zTp6bhVaC641jd9tY0TRP5bJ8oEyxRfFB7SsfapStQMd2vl+uaQPmp2ECt1x
YxUNmWaqFvt0mDzishRMsREUyDGBXpz35ulrZgsvVQ36fZEoiUZxSeimcwNHwuc35MtELbx0DfOw
8YiVtHcn1Wbi2ee2sC5w3/94tHlMFjHNJKaihsLVlasOINGJHO2iMWQo8n0Xq8FEVClk7BT8jeik
NoCCtSLYUyMRgahCKEtcfH3RdtOc1dJ4xjWV00JwR7qA97mu02yv+ntf2cAZ+THE/cCjFjde2kOj
exXpJd8Pnk6RzwhU/Xb4IxpIYKdli7Z+HPkoCu/W/KbqBdoYExU8vMXCNRGHISCr/p5B7ZWNB4/i
c49jTTSr46Iyze5Ny3/vEE0rDgYetC07EEmNa5nhMS7yGyIszhgZt4faHrFeUc0m7EtXCHftW123
52yUawinBiCPPjepuiuzl+yU3HcsGy9AFJvci4pEromm1GWLmOn+I+IaaG4quBflq1QevzUkj8C3
znHyYCQjszQ41cYrpdrUxZFFeqsufIK2XWJaZupISLKNokPetS/HW1Up5OHpmvDLTiHCc1F8Vs3f
0OnN8x3Q3hP9J/gvyEnAjnV9EM0qfCvvE9LPS2MA4+Pwg/e4ykBp8JcPXMuWnSRWvOoXodr4ZX9L
rn+x1VaD+zQJmssjyTkH6+w7DnUp+KAcrDqtzSSEOuI8KD0Cy36IBOd4rL4n4XjymL3QOgKR0q2X
Ck4QJsVTTcESkVwTXkVrM/XdZnynV6iB6NAS59U++tF0Sy7z813l0/5a/OTv0yh/encZJg/oUKZQ
wv0oxgl6c3pF1clC9OsPf6DSfXxug31FKwcNcFsCjDItTI5fqnZktt9GBV+Z8dV0YEXhCG2WQ8TG
Qp2ZJJnBJApJD91Z7jlAWLXmFPVKs3GoWjJLhIcBTWOVZ6/XUV7EltPh1H86sdS/9sCKpX9rnaTS
oEFOAs7TeTtZKi65tIPTIHvvqy5MrHc7Eu/haWlzXqdllgOM+J56DURHsR1MfnEaVbz4AbnnT62Z
iV1AYV3fEGSs9qw4DKoRZLG4TV/xDe8za3FoXCL0FZXIM9dWr74HVtQeVVgv4TjtITOr16Mwafgd
8bxK9wWjHZPJK2SWuKCH/CHx9RGOM0HoCqkJPurgE/KNcl43yNYOaX1e8AEVPieeXUWzazoYvDmN
YpHCqHuh4p5XntIY45uQxJNKEWNQIRNIW4o+4VqaKo4KbVMa95IVbHUDC9TNLcueM5F58FZLxnHO
pMPgt7en0alj7s2mRAId3T1e/7TiYzhmvtW7rPagPI3MTavMGDw3s6A5Zlxf6+rwJbbCeMx3qseD
a6DoZRDKijrYT4UdIJO6uAOVrRoI6M14l5IJ3aEs0InYCK4eTe/TqNLj4pPbWQy1FwDpCvi4Hljm
BYM20BpiqCbSAErBNyj6BFJVkGKwSegJEEtjM5FY4UTZIF4bMOB7nWjcaONXN9JLiVab/VVhL0Tb
sxKwn6bTSBcVmW0ZRLhQmQ0dcy59QuyA1uxFZ4dnHzLGbqTF3neBCJ8rEQkaqacSlH8kRceT+ptL
d90Ylz5h4Z8kHibVcKPDlv0ypgRUlVoNXZZQu5LdcKYwMKbSrqwPhqUCeiICjWAWd1E/FEhVOL6d
m1+E6d9xqHgUedWFDdR+ZaCpzDS5P0xyKuYqKKlTvUY75i8t3UisXg/eLsyF0GEw3dv/D4eymLdB
CKOrw0TMR+LDDVpfjOaQkZoc4gwUFjSZuNRYJDAkb0LBzY32THJ+vsNSWdqakFHeXvP2WOMSRnHB
W3JReX7Gqw+PsEtSXcQQ7wu6YX1ivSdVKWdB5tv1JxAOuqXEWhuvd/XGCFSMvJhTGHOO801GYDJV
5jcTlhf+RT0+NxhvrORFXkjTynu8gnsGYQ1XYUSqybg7TiNg5E4VdAhtyRaCJ9eQEexyXzwHg/xl
WXbaYew1PDVOmGSmHW2pr16uDiQGjzCuQ7LJils0MMvjxUEaKsWLW1ioJukv9+C8XKwKOUsxlZ2G
pHiwH+aTF2+TBcE7v1undzxtt6VEAswLv0/9O4Ds65qZwxI9Pg3SgzTFHNcMF5BPfKv2uyE0GuFz
xMBeKqMJCtyOjjYY1fpMrfdEwYZ8f5ZU+BkXu9UdQYwbG2Zl/rstltykI8P2DtFYObKEgjU4gymc
MnNNrfqYe4nK5qxCpF1Fb0sgnCXyKTYLMxpipLnE78XWVm+9V+0MFwY9fg0hhSgqQVmsm1Rp3C0L
ai3h9DGgZXLQE3c1XqG32cGHxaQWuPwg2GDTaL/siT5KE0YeHmZ2/Y45/AIrYKBmFnLNGH0HLp+u
Db5z09vXlxLMp4ghZTtmQ9cqcqHc2mrkupLqpNJd6rrFMQtENT0wWKwNE7Ulw4m8+Q3QFqnpFF2q
7tQ+1/cfxYQxdiF0ZLrU9zCctB6udvpkme4XOZ7v3rckExEtL9f1ejhTzkqjfgEq8SPCsfrPaU2d
ePPO35We8p/OuzO2X/rb37Gb5Mw6TeLmOTOvhFQojuop2lqOevyLQcdnEFm5dKHWUvpKjSg6YNz4
ZFPNYamPuEfyanIVq73GOyj2PVXlZtBkZDX0qolRanFUERH9ZlBzVTagCrBwbmFjbgW9OefvMbqr
yMT3DLCxj/pN1ZGZ1HkJNPqCbLrhsC5Jl2lsZyYPkeBmUVU5qORWlRSpr89zG3/Cq3rR6RF8Bxt7
Hazrpg6F7GCZEPcrfDF1myv/jrE6+KhJontPZ/atuL/UTC1T49SGLhUxnGBgaFmOCsGp5CnMBgh6
Udivd7ULGl9+tZBkKbriq+J4tUZEeBev0BZePqXKO9r6C898golFYpkF+KDmkc7I8LTfdM0jjYMm
gnXEhDIypqNgfVQp4/2YQ0pMnFnAA1jQtc2ENj4x9odCPP4KZ8DGLiiaD8b6Kygasc1NJqN+M//M
kcD7RUaNwBZH40KQLKdDmHpxfJV7mjZpBG4XWsJyLzqy3O4lrrgZPY2u6ooRwiIe8ut59yYL7E58
IATvN7Krr1m3ioZN8vWOMeXWwudgYIDF5z+FsW/jQe1V2FHOuVahg2mPeZOWrONhX/GfICOs/XQR
0LUye+h10hHKzPBOUMwF34d3ZkhG9WrO/bdJdWt3HwNd9uBjfSQM7bWykDyju4V5j6wW6/X7YEqC
/MDe20bBTTfba2AN6LcjWceZDNfSRgD2hE+Uv+efUjnKKte7zMRcR4tzSYPz2m4pm+uQMPxKOj1u
XHwGkrEmkqACfdMu6Qe3vHLxPjZG8gb9QmPRsb2V1wu9xIKusiU9fNJYM22OCT1JSeYpPpwE3CYW
VVkucfvxRBvrTAggVsyUePdh+4Y0scXFDZMjGCtzOIjusXj1UtQ5eTyKtRFWfd0aWBrbn8AO4you
ot7kBAYmQybGCuw+0EryqQo1QmMX94kp0GyBcCuvSzlq3c7GqUu0jgKD7y0n6X41IZO+19Gt5HYZ
jK16IiQmQasuAgvEIpEnrW2i9KwAsNNaPJiwJUsxnI6IoeouIZfJZ+cehWRAGkmE8MEQRq/1kNgb
AGzgcjYG1lITz0WsPj1bMiuVEhwkvZwXeJ+WsfQ7X8K2hbCzRPlvKzoTqMNp1lSL+/+8gVb2OleS
qMVWwm/vl6BtBCDdVGuf75iNuNOnUatKbIn63wTebSffrKHRSkud/G+WYV047tuI9ljx/3u1jCNP
RP+r+OLeKJUMa38uf1QkbyA8nkHfRuL1vQdnvW8n9gTULos8rfevaIZIh5QRKbWoixyfKz5qXAt5
WIrIOyoXkMVwraEVpJdyZcAFIwHQ/u0a88wM8fMVXU5t6POLNxpeFzEzsT/vP/Gd1Qn5Y859laMG
qstIRxiOz6mNOiTG5vDvNDeA68KLJVoELHS9BZMJ70aPNla2Nz0qfWp+Zk3gEusbP0Rea0HnEZqj
ZcF681T77NjZypg55EBZH6luMjQgLuA0NqBat5s4+0CnbgmCREp6GsQY2PYHwKwXeILTOPiTtYzd
9vRfyp3X8r5HyM88a75/5CywtSp2BKsYDnSKo9kGcN5VBsbleoJnHjSi7xO3yXMYYT1zlm4QZ1df
UqhbVaWOtgteMP2eW4a57QB/vvWDBE066ANnNjfTaB6Xjvhqq7i1KQsjzElt4p01sb0WVp/4u3Rt
evM1E9zwf4KyPsmHX7M6Z4FoznoS1QMUW6WcdlAT50Dnq9rVqROvvqkpuYUwm2oiLaZAE1Q4/u8k
XPNlbe8A+sg0euDROlFdl/A+EiTA+UgZpR8zipGqZxUdAc9aPJ4vGauhuhnVzIGFBe8cbIwCuZF0
QS4HM87qqM9YbJJ1GveZ9NmT30QOhImGkzU59rm4GD8Fqc1kVnfcTOOmvXmAralv720IMmUC5hhT
RHrnpfUFGmwv/dOaLiv0ggt1YjNE++/EiM+P1iovLPptm2QyGzeGBEDlxOyYpTXgMCedzk/9ZHl0
bWLjFlEvVChqxxGGwJNKy+5sq9627flNiNdiJMLbRuqSf4wB1gqP9clIGMDraVOZCTr1wenZSJyU
MXo4FTCceMBh/0biw+7eHSxAA5RqxXfj06MZAISYQyQ85KJJ450paRtBlHrCqiThstYr/oMtKpuq
JA69De/dF1UQd/oV1xloA1FSulmKbICJ/6eVXqBsp8bol33RHvOnhxn5AeBMKuCjPp92r9JJCSvc
7ivMiswo1aBSQEsDQHzoBKLNFjJIssosvPG3oonX2TeXklzY7NMLZ2vcKdTnGx0grBtUfz80jGXJ
4IjtMSMtaMosx4KeZm4YdcKLCq5H0ecuddfze4QK3YJnLn1aFaUarPknLiAhBOzTZJmWpovnmOqT
oGvbK/3BSipdvODu1mP+Id0pV5zwvb9alrI5HnKFcaVc8fObaIG8oNfMGfNG0M8vHGKfROyucYFH
zHHevU/NXD8Zdtkm2oE6M/TI8cLq1Y81fJaQlApWysqOcQH6H+93oQ7Okr8Lj4NTBw6XeyTqA/or
bEM+ka5vKJVh/t0lzzPeYSRXsfeM+BlGmJKT9h9xVeohpXuMHwTYuJR5p7AvnDYLLsNiXGZZmbQf
yxGBiito9eJ4CjM4wGOexyc9tDB/U1XQQtFbdBysxHBg/RWGAkMZO/l4MC8lbX4qdb3hjOIQInCM
9GYuAh+96w7wVH8YYZ6Txy+0/rpCdlOHZ3WYrE5hM/qUln1QW9SzTBY9PMQz2w7mbOu3iGb5bhcP
pBDyCuLeKhTvZEqIukbMKBkhss5sn27bexjWgIlQfA3z7257zahocX2rC1KIfdrqAC0m8B5RTMx8
Q9neJASbTwJF5LK/TI1PDZCJJfUCeLLAbBuDF7XdQcUX/JpxI6ALt14xcysG6iigov0ikfgL3PiO
28hE7a+Oeibqb7vrzupiitL9kqVUN/JY71BeGudr9qZjRWCB6CQoeqiUsH7w4yNQuyXqn/Ta0vje
UOEW437GvaOLc7ugZrCQQXNa6zjYsLXelvneWe4UmZYXc2c5GFnInq3Zso1CbZ0buPzR7Zkv/djg
gNk1QLH+bohHZutgYei55JbLFGL5JH+z1GA01cKztPfaZCrX8Sm+KN+g2xidIQveeGKVwrtqllgr
GZgwEZ553Io5/+DTtEoxXIkJmsnEvdZUSNKSD5GtQxEne8LqUFo4u6ywyVEUhyh4Dan76F4/BhSA
ZWKIw4pqWnrz2nDURcqohzRFAdGH13yQiVA0BQh+mK+Qr6Yl+g7GXQxHkH8XXu3RUWH2xjNn+Y+C
BNLuHxaFbNinA2BzdRpIPHQ0NuQDthgB3qKLZEqF0eDXCVotPm1aWD7l7FR2hmrr8pkUQBflLOq6
6+f1X2hGbO00NRluvSIVOcuPAu9hopqCynkRhckcTeD7mTCfH/0Whc2jMqycmmoDibe6M/htrgE/
5gdewqvGWE3js9+G4TRyfCivfFqKMcQOXBe7mcE67HMajcDDLN5DB9N26AN8Ha7kuxPyG8m/iqE2
7Z8nZc1AYMFZU4ob1wEXwGwcbuZNIrLhJ3Z3kpk7nBX/vC3SfEMXQWD6J2eOVFYX7YUphoWDaqh+
nWRwWytWyvbaO5Nb1xaMe8BJJPxO8RVvSRYMinCBqvWnEoCwRdDRsNQOCLNk0sCRWOrM0zmz2kOT
7INtWFz+73S3cUgEzJ+eEh1com8FYHWGNnLmIDVV7Y65sVtQGOcS+mfqIGYcx1K4jBEPB3V68Gpp
AQS6PEJ5X5cKFVg86ccLZEMc060ixVE1hvjOqd0GK7LFHz7uehBqcKE2uLsbHIwSZLbUCVZzy15O
NYiatscmXs9AAGIEkDe1QVUYi4dNdSYh4n+dvzP+1h7Q679x24eOWkmO8C1wyzCjzVhqvgG/58Z0
xLoFb/UktHcigjgGLCoEB49rh/xoHvOFBk8MxRluw6lqfYiIHO18ZGTaVR1xiXakJuBqHHSzqqix
0uRcd67AGNk2G2xW+R/wWnJ/cRPA6tQsZw32zffgIixyk0mIu8HKfr4Z94LGIqWVoVt0yB7HCSqs
ywXpIpHksiP69wf0bW0IpprHxlSTmrJPVWb8kMsrqO8noV5ww2eo59sefCepj7woASsvk4gXly/y
4YJvkFQ+2wItXtsgc8+HTlrXYcWqPWJR6r0ElnWfAG3TAKBuXIO5Vi08NkdIIOim1YRUgj20ezzA
KtCWUEFk1vUIQ69x6I95B1Y5pl5EvOb/nVhwp7YpOp5UFpkWfMS+ShLV5wnrwZgMHuA25Y3d/aNy
8IB6ZjceSGTwdMvTawNYUo1+idzRRu5rFbHdP83Aukv3jloWumskt/CNw0eMDsba5y5QNHE7xzDy
bAWC2Ui2i17/YQGfUPEVIBLPtVwEcMvWVrTif/QWtjUsa/tVjregQK7fGPsOBXzRnfE5WK6JUDfu
5G8Gily9BliPHm6VRAIHeQKgKu0OydXqp5JpitjuESgvv1fTg6IQWQrlguc7I8cX1ri1Fjdxtfjc
Os/tvnGTqyZU+nimia5lYcjrEGZL8AhK5cbWmGbFnaYuq3Qq2GdWV4v0hPZkdlw2Q8BIO2qcI4wQ
WSBpAXfzVcrAxb+AVx2/5Mxc3OBh2rqQgiTq8FWpmQ+5rkxXkOHZI/pRTrruXlOOyXQ4IxbAoKOz
lifS6XlXP2IMScnJkyOzsmp5U4cc7EGQlPWui3vgodcuQ2LSTtZgyQF5viO4YwX5lg8Wk/TJhtfj
bJbwt5Sb58AHaYtu/gAd1eq1AnxceVbWzRni2k5oVGXop0R4WMlqWOmRR70l+RcU54r1cRFu622W
WZVqQw1k3N3ViFjtkP+/FWTwuTP/UdEcgq81wyAH3zo5/zsR0UDQ+YIKO+IQ4qETtKYzP6fs1hYt
XPesZoOMC7bQTRKbal+5eEgU/EIA5TZlx1f/SU48s90zJ6Gkbte8iGpgrcvoGVpRwnMsQlUVSoOL
p73Y0zjEjtO6cr/33rTQ+Q+KB0twTa9rhs3wdHu2lNXvLpSDWpaIFGaNEDFl43SQ14PcWVl/MZl7
9AN+iCkvjfn55J2UwXCJZae+UoVl0bW25ftZ2I34JXKj0D0gq5tF2y6ukArbIJI5o4QQvu5XKjtX
00V04xNiM7fZ83wg4qjWJQjhwgogP5O7TQ+97WqP1/svmg3QibBA3qoF7PRTlssT9Q4QaV3wLf9J
nQeRcMQQyYEbjh+iCBpNL+oE3OYs5/zMeVhfdx7bcq4jrKza/3HT76YsAEUc6e8cpFFlzEOepQ8D
ssoazDY+0u0LHUL+PO19y+DKZ8WeDXebJfUprwfLfvTxNMpyrapu42qsoDL7lsMB5LQbVPzzI3pp
Tw2+LpZvQi2nGPjJGo8vqoP5IRR4DKGRx3eCj3ebH303hcaN6BStFh1yzaVxG3FZoz+omDQi4pH4
+jZh3o9oUXC+7GXZziBVbnu4ux1xXE/SWQ84x1kLTGike5Tvncz0pfrKsMWpCjIO7cQXXp5VsTQV
f5dW3xaY9YJJ3aFA6q49CIW8q7f7oIpig1K5scWQG5rN8M/ImUB4jIcCYmHTDyfS6W7m6bvIR74b
YiH07UVlz8gZRMPd0dHyOENVExMr3wMjOvmY/T+ZGjnpyCVr5QVh/Oax3xVZCegwzbKWJmUYRrcC
luS8MWnq29BWqSQc/EBCFjkMjvo+gXpGsHn8Xa4htkK1N/EL4Sd6txxewhoN+hrp2wZe4B3ahA2J
Ph+nkRDlM5hw+ogWYl5v9KP5eP3OZxigJ+HfWNwxQfLks1GOEYW2zNhWCyz3JaPytQ9J2z6Wlf5Z
9v+6NxADfp8P08eX+1OUyUX5CcULLvdLEpQkwQp/dOotHRvF5P/7uIvKzxVqr6LtdXVSn+T7T8BF
FNOy5bZnI668jFgGywzBADspPxDC9mst4FxgpESRcAwF53bRYha6CtvDoOAZeE5no0RhlJUYjKz1
NCiQJfaBzKCLtbPLiTHeOoc6tDrxn5v9GBkdInaE7S1xK/X4+PHWkK9v7dTi5Ra0chcBMgnpKrLb
9iQduHubR/SayfNqcF9PnhmNmNhxnnzzI/PNz7BfNdGtuQTgXXOy0/YHPDKUaOlYRt7DCF7HohIJ
GSh9nixxo0mAdHqbR70NZJFJPArlNJWPPMC15CTmIoqQAp4Ua5Ttg1nDPwXiwOagu68tRTiZ8jE6
Yqny8nIVFP8oTKrSUn6xX9+PG6aNDiJ1W0XDco9tDNqjezSVu/uIf2LxCVDFs1AJXLIicsl/1GSA
MRpP1wn078ukZVKOkiV9tjzxbSwhfbitDPBukm+VatxjQ5UKK3g9zFvyHPt1F7RICT3P5PGCYtJg
hnsyRPTc+/k05lL90KXSouJnpTgGO+umRZU9/uN/ifGCmJTRoWBoRUZhw8nw8naF8uC8IdAzoaVB
axo5S1gLzTGy5VJSbmjOCtcO8Lm7yy3qbJG21REaYTFGpWrHrubDGDmuTg3RxaG8o/M4JBqWA4ZY
XHIl+MpwqtcCIW1EmGyc37UibtqLuEJXqzMRR0Tj/Dk4qB7hDH/FCHi1vAccBiRoYjc3YJKd78q1
8rSFPJlTZS/Xn0IJZ4ERMNv7MpJEbUzB+0PL1j+oWuM23ALRcSGXFmgr2QpvLSM6IM/VM6J+j01P
EG7U0bB3nKo4fyGLLdkbfAiZK6ftQ0sTg9YEbmG7tLQ9UhyppvI0+HunmtuRQme5kGofJ2fuzG3u
u7rVA0Gm+2TjeJxgu/8GBntgiQLQ4dGb0trf3N0ikYRyXZ58n3Pri1gASoiyyd3LM0TQUkfGCQat
0K1K1GEhoAvtK1oRgGmPeV3Vg2wecgbzvIdVMQ8i4BrtheFwgQuUlQiopiQnLHgT+x3wfhIeM/th
v/boOKQeIEl+Q2txNqUVobrMDc6c0S4mStL9fpEETiqL9iGXEriVrjcgTiAWqVyqmx6iuRK3gEsP
wIfM0thYCQbadCEyOI4fi9vulBPsCMXPCOybl9Esl5UfAIGST1sCFlChNzwlmoWSOb+kp3jNog8G
/uVMXPS+atRLfjiPRt5NCHkM/9KhyLRsBlgdy3dtdir03NVbm77WTz4zGRbb1sKgm+0zo7G/D+Df
dOAjSgRL5CkNB4MEjqO193V+uqygjZyIV5IMuCxvbIJH+JxPeDA1PqhL9nXKp5pZq7pHteB/9Giy
F/PA+qYyAUZUp92FKWL89ymevXiYtY4h+7voSazk67PMGccs2Fs5XjGjEg/KCPzDMDp+cLD+IhRo
/fDFzZrFd7jfHXljb7hdCZAE12VMLXjfeOjobfzmSjVWaVISyNjigLDrEKUk5BQ7MvTHMhv9i/gZ
MHHk48DYZTpVrMMeZM3M7A60lHQrojaBNsBWf5xmihPBZ59fXKEmPeQN2LuohWIZlK/e9bw6lh5e
OzYjTha2us5PrIjqRrZP9HLd0+3Fvb5IcJqw2LfEajsEXOSbRN6qmhFZX1s+AauU6Rf2MlK6nikH
wn6ajRoObKA+FH7jfLqEwkgDI9u17SNTLI1czgOVNaABdKltYIAj7o01S6PL/mO5e+taO9NMM+Ob
gq7OIzkZAmG7XWJNnltKZOXd62uodoRxS5O0SUiLlmMwPKIt2BO2YhOidNidFM1xbELDraM1Valn
TrHJ4bunqBJV0RVO55/1VvPwA3px2nBhI1ZWUREnnaNVfKYZrbCvvKOzOEg8JusQN/eWdJBHB5Oh
1VHixHJXRMHzmYWsYk9M5WS2ZEtVvaQ2SxlEZT8Uy2ZKk8dnn/GfTkIKmCUSfvKNHedOIdNakZKN
0HL3WfAFacVk/8V/1F+u9OrmvpJHQ+1Byo+cBcKJAFn5BoeUT48egInFI5QddwT1xfiSxPDA6Miw
29aW9lr8nZJ6U38UcXmN3l87hGbnvCueIbGW3m+pVtCD3bk32yhH0ifeIhXliVCUXIceruymz/w4
0bSNTVSvVSjOnm9RMt+4NBf1414xYlTIOBB/2h5lUwbMYIKgbogzg61wmjX/lp11qmUvrpZN4NJS
gwyQNcO9qWIXERODn6XQXjD0NqoWEubWP9APmdDydrg/bgNNybpAbfFGLJWrcDbAjQ1ZpfuQ8NPs
MeW6saT7RFp5jSnnjJTE6SH5BQ/d3/WajL0z9hvG/7PyDT/ZHgStLCAXp4IjtsHqAQVZvXC5tGiy
EKdqCx+3lc+usxC5kFr11Xq0QQPz6X84Iwv1VNvR4F5QG5taMgrEPiVv3kAQ2vX+twglSlT9fxdB
J8SL5aSsOJLEIRom0KAuDD833zHQqEjqlkfiMGAuQC61RT+mYuL/3yptEJzXimKG6d4hQzpPf8Mm
lZY4JdD+WmoHAjzLroWnX9/915fkASsUxuzlEFOJLYv59zljRBl5u02bmRBHzZIkMv1QayqkYQev
AfstDqzIOHVPUG4ZDsNOwtRlkRML00sMUC/MGpJTteaC0mR5U7g6QfMzYe+XN3bPs8vzkZbInq5q
j9nKPPakj/eqHRHh7zRA/Bqwj4FeuYj48RSk8pcixtoEVY+O64pzSW0PabEMdzi64++iZv7PjZBb
V39FhsQiqBAzC1cUOyh5cUeeaE/TnkHegTtMn+Ek/iVJ+K1P/p1mxONdO8XcAHoNAMqC7vzMe+ur
NgYWNW3G5Wil1CkTUBR5DwzVwU1wFc++tFY7fQ/7YMKjgIHsTamEDCE4OVk8WSIJTBiSYuVK5zBm
1QUOBc8Xxx0aO1L/ZYJ7QuYXdT9NTwMZa4l+v1bHknhHBb1+ycZQG/S7RQjFAnDGYLJn0OkBMuLG
jOAGMRghrH848yufjrA7y030rQFFER/WPK/RnfSd4KDSXGmp8wC4KvNIXeQ0QsNCfKCLpp6qTnlm
ZljS3K5f/2cN/OXzpP6Iy2A/WPvzTnpA/5RDrxnDNakw7pHptYNuK4/c7Vacxx/xU1hIqxzQO8jJ
62M4yVFXY+Z4T/Gy75ZPoNBIobLrgZhc7JAkd5MJuTfueCd19naRh+nLFHlIVxmJNOlskvWXKn4p
SRgxGdqBh2mbc50dJzQ978ASlw5wKF+Ivxgs9rEO3ZFWxURgdfb/fxMa6M6AS+1Akre1Y4lSPczl
EcZ2XECcScdwzIOHkTlwq3xgF6Uq/TkaGwYa3gvfNZTkqT0VdGbhIeNCWmh7nm2EAqVFJB7gJhcz
2skq3Tg/c6eC2zdYGI7cs1nwqaNGkmzxYbjF2m+iB0PXkEShjj+IpoVg6IzI/v3ixNci13YsdeIe
cfpfqz6d15bbKtdjBOtSK6QnlhrzdmFDLilizAgZmc9V+K8KzqqPMjMd7puoRBYumJ6ib1iC2GW6
8QY7yDYO0O61a5/34McNruyUX8vdlWxS8ArktwpHqkHMAiDljUzNFkt2nsIiubTw9g4I4ZhDnxRA
Ivd5JhewIKItWCWsxQhL5QFq82kMnwlNYxwLgnqdGdpEravPNGYYuqTDglsMOPyYXr37TUB7C7CG
QB3dK3KZf/Rp2IFTZ8kyYtdduc4ue4n2PEtiDC7XDGt0Ja+X+GEhSK0iFVmTNy1tknujqWeVh4uO
zM7F2zyU6uQ0XRYl6ae6yQE9i/qA17tFqG0GEvuCPtJZ32jbftGzHbunwA3HfUb13V2bEUdLZsb/
PSz2fzdD4q1VFMltxkJytWu5djty/fbNy+gA/5tMMQqYWFPZIJutfec1OqDoYCX0B2guw3IpENnO
Enbyr3GYZGaaU7iPxIxluPOV8kdJefQsGBkz2bPc8pin1MrtxcW+UzsGY7nMByZT00b8c5LebDuj
eIy2ZtO6Gx9JdZiJPpl/V7pGLmhd6/ktOQZp2TNioZVKQTGBR6y+GMsFX5AZiwKFxKCEJkcB2oV/
X4/d1WH1Kq5FUGVvMyEy5V6LHsTQAu3XNBlqBwqoLTHjJkk0TfYliwhlS1/3E8JPHqx+MW0jaVsq
vL6gg3pwdB6Xp8CyiCljSBR0xngMO0x0Z8LwgvEyuGRN+xyHux0V4hEhwsgpj4qXBcEghHf6PJwF
NpyP7cW7zY/3H6PDoEuuwQ5xosx2PrqzNT9pPT8Nz+oSk9zXkDcEfPQbFz9ehGliXUkT6jNFWLhu
yG7tSdUmtxz3uqi44TLqPo1CVDxy9uoWJZJMKvRQRZAnWXToJtXVzmYAzsx9b6vX8h92Wde4UUDf
Gc47jikPg/xGUYxX+7zVI9N6C5wj85HrtQHvJwrEoz5aIAVHQP+jMFOU4Q6LV+WOLiazLl1adY2i
yNDnKnHiyVqYkZD4c0y7oZDZkpq5tEETnVkVqCYkR85xdIDG6ZJiONO/CHShSZA9P51wu5ZAmkr4
WKBDYLehjL2CwwLU5uAbladZZI7NaAvISw4kPU0icriuBmFPhKzGoq6a00KhA0COhoaSTrKWl1YH
Gi57cP5CUKRESHgfuikYb6xi6qElJ8gC1bL24MdJ6vmfbp8FxZIuFjfoqq3LcP0yV1dOr9vtPM9/
okTdw+HY2uKG2hcy7g0KVol/OskiffrpT5h07OnVdSdxDtkDSu+YI6Rgw0AuJaNsIMKNfiUCHlAE
bG1F40IlPM9fWGFFUesMi1lngyMOBykEt0eixuGwS9ATTWTK92Y6qfNlAHdJuQAnD0XFEnLl1fU0
B6Iz++PWr2IDeeN+rMhJ1rgHqCM8/YJVD2vgp0agKmvp5kPDSNEH3WKJmxZRUf/L0UiX4JoxVYYG
XksMpTKTcqENb7Uvv/6A04jJqUZbxgENMkNjzEfsGm9oCKs5WwRh5sxRFc4V8wrsaeGf/Iq0Vh0H
QZtXMEFuLBqFalSXY0SX9/vLEQleptuj8/cJgmmPigjbmjj5UXTLyfNnyJvWXXUQqSpUl2rvmkv0
II6kYDrLsaBtgPGj0tgH4tw3HnBSHO2E0VYnreNSvZ2FFPhcly/BrPQR8NB7fCrn5SG+uGF5fefA
Oz+MYGGpZ9VI6oWPN9pxS2uh+pElr1fUHVe0BXkfJtmUXJTMThvR1F/Qoaedz+5kF4xYNlOPpVig
WQBOXgp/Pma4UpnurnuuDHLNGv1r57Ehb0iadQOW4d+zyktPbfIh4hNco2/CgkViv3D8JbKhGm38
n4nkwA+UbF+Om1pdG7R2kloxVoK9+94l4yUTzxWsFTwAreNlbVO5QYqFFA/QelVXXxaLma3UAnLz
7EcoxCaBx5sVnsJ7Mgp5Np7PrMiInaUWi+Azbl6j2VZ7A5UOZ6o0PwlU6wITd8U79pk/s+ftRd21
XuCPX+ZGlORJshSm3+GzuobGIQURko0+0ESpJCMvl4P+Ijsw9cA+I1ZB4/sqC3WPpNbvVnf4iYeE
6SPZ2DA0GiZ8mo6th1iiH+/Gs5YLT2A4Bx09Y5fyTFUgKfh+ifh/QhtqZofuaAzhdNvES1R+BiCq
U9i5cD0Gm6Nm0U+APMEquxOdUqm5+XXJ2ciBzwurWqQTqarW2TJ4ZOvs0eIRsI1VFOMMNPiLOH+N
RC/jtHkL+8i15bP+FzeJ28n6foGWJd1rnoY01hhNY7fPYcZvJN7jYSTl4whSu2LfvO/QwecjVZgB
dF9vwdVebHBNfUSaVqHDiPZdbncWOTXCatCjZ1pL8jL9YcIy6y4psbSvtBByK/s5AnJ9srtVFOnq
WZfjWLfaEhdMqHTvuWiCFXuWR6x2Z+kRbRnL2uNpsWEiXuMWNCumSdcdggTZCse+HLWSnkgmLnyS
/wobUUkI6K6QdVenYhI8rPiTujVxLORDpzHlG0W7nqM9U3ev5gG+hvO84WYzSL370ES4oquw8ytf
3BZBmCxxC6KFNVgMoOVFn6Y/X3LmuQCXsIk1QrtFvx47Gnm8gCFLVI2kVwmcXZUoVWy326ccUB55
RikPcyg6EfF4f1VJzpg0ziUiGoCXM21q/zWjcLA9jR7uUR2hAN4FQzR3F5eeAoCyZWRTWimwvyuO
LJCZzd7y2jNmKvRVTVyh5eQuC35TLLa/KbNfRNDq0vTL7wEAYpup+4JJsabm8QFQbI3C4QP7vCJ3
Iubwp/W6tR+batTdd4uFpPEqydsBgAhWrIy2ktDIlOxzAjoned9FR6w5x8Gi6/HlBtAaWT2aL+5e
ctABqi/nfnmfmc81YvIbfcRCrGez44fd7mn9tTAauvggAzZnyvOI6KRV3+iTZIzjubF0OWbaa2q3
3TcvyJakGqEi9UNeyH7ewGhzY3VBCml1ekyYdNuIyfB1WDzmrVWX8KrgbP/kFFanlOG0wsrUyBta
ttKLsyTD4eDKj8rvJoBWkts89p2q6TiBauDPzEUX0Zpn4ckIwM0SezO9ksGdFoWkcGgGNSq3ouOE
7PuJtQFjIS/vg5WKjWeKrQw4Cmt4RFVoE0N9ui05hhKcFMr6qHiHug+I4wLegcBHhaBdTVrEmZr+
XV4D/iqZQOh5JE9MSWZlgPlu5HRWnpRd59lOUNxZUy5YzcIXBmWkLARoh50nYsoCQCCsuA2RjR7V
jImZGQLltjP/80WIOB6ZtAZLKhAxWg+ba5lKIBaCRHzLQEyNyq2C43O61jTinOtIl7l9dMCjAYCe
lAaNXDyG4qpZVIc0/glV6XEDOMPl4gz/Vdj2NRXRnJNEugtVmkBnHzkz4INCX2JbpLGbc9YnzAsD
H6pggDiAUc0eIn9T7e8JelBp6Q+e9LZes/8JxMBbkp9iNZ1Ee+FuFDAQwo90UULxElePrmc2Y50i
9L59rTaIocVspnrPw0TX9h3CL9iaTLDXmj4b+UDEI32n5lMaaZE/5x316lacPJq1pN1kqBGfZny0
FhXjPZFm6xkhdCkDYYJE+Q768Scg8Af9PkTTd2WTjA5rLIvx/ZHCcNOBURziDA++Hxvr4mHyv6ju
elY3GirZX/Qmil5wrIDxKLmcqraRISKrkxZK+ZHqYXlu+7GWxwuU4VSe+pl/zL7cCfNomY7zUGZR
cqK02nAo4kgTaJAMRpKZB9iNxw1RBwbRJa/WZQd2q3Rn1//JrctwssA1NRSdcz1+muTfdC39tVcK
6PVKzofATG5/Xl1BTYjQ1p6CF1EpDpidjKLI9zJDyoGrnZL2M3TAu1kEvwmhS+VfOY8W8AaClTfZ
05xlXC9LYF2EQG459rqsB6vHqD+QH3r54gYrTVuPS0peqstrRZB3BtjyUk/7lApeDF3bEZQwL5Sq
5ebSRLocjiAvnXe1myvbzOC6NDcqRGi3IXp6FLe16tRJVIaZvZcGqLgI1DPt5b1+Bd29ZBErs2+g
vwmcAyP24cJjNMHImWx+E6AaIQXvslOCfnMYSiSYUz92KnHh7jpnjXwQXKDpWIs8QUp5+wPMgD2W
hwqFj1OCgDH45uEqFeRyygT1+5297/GboyCdkb+aaTWKoBYzaDLXYRLsy4QqSimre8kkQRgCWbFx
PgRczi0F9qTSGcbaLQWgKHmDU37bbymSWiuk4jFjQXWVWovQc6+a/+p8jWd+nbKJZYIHTJE2xcPF
8rBVB2Onps1i/UpRtH/55cs8BcxWn5qMwhqG0dNqS2HPSY4rrVaWf/wnr+eRI0656BnWTPZUYHgb
BExhgSzjh3PR7qhCXGgDjJWb0ifr4/TmTWGAiWmv7rRaOuisFJFTmeCstf0EWN/DmqfEyccw1b7R
qo0V98ioQhUYNSzY4ovfZqiEmd75Pimc2W5sjLq3pO4soNnF3sJbK2RN1+/ycZ4TPZ+S8/Al5qQD
fP71dWKy6HR6J2GRVVRvCCkAk+OFJM9J8R9yp7nETsIxIhoLpTfPlNmQ4F7Hl9VqtQwFh++68amD
9XYWu6uvXSpVLbc1I3v0djWt+g+K4WQyMRR6Q3BLFpAApSWoOUrZG+3uGq/29gd0OZUHWe1VCzQh
RhGaBKosigCAYwD0q92HDa9KZ6VAiu9lbOc9rbeQlR6rnF6TdEGB1wq0LIahowS3w1KtX935sfDy
aoZb1DpbK2NHi40KwYPNJuj6G0/KjQSAOLjfFSa3EKLUI1O8AF619NgFSl5/fdLPjX4iwOYBbKcN
UtkYeJ+mor7NuZGT0pRqeVFKvwR2yVQgSt5cptE4HV+sG3xqwn2iWAW7Es5NbYdTvL7WHoXcIQx8
hHBfl7kdtTtVqieMZh7GFe+MVs4tp2IIGeJaujJKuQrSq975gLOXWEXu1mhTiZjO3biQKtyTDgDB
JynxcXovwI7i0tsDmug4Bzty8AmaNwDcc+pZ4PKmcgU9Frm5mca7PDZEiZd9XOOuTxWKg/jCjKMt
P4w2vQGJ6dnZx9XdwRW84c0xEdBLf53EANswnNUWSlPAZaKW/YNF+TXzTR7VHFWj6cxL6dgxrnLv
NFR/BjMCtK4ww8/f3v+z3d80TZxOfVr5Xmiytcc+9kfKC666X8lRj7RTOpWVsk1/0+jK7S+qcIWC
GHu9F0/lfOEO1NggR3M3pqMES8c/KF3v+3rS99JaHeglu0fhiHMHIJ4ACIWLZSf5WAHZhq/vVt+P
IfQNFH03l6cN1mSVN1ckT00K/wtBALEttW8OSYAm6ne/d0wQHx1RWCx9f83WckynO8iFnWmioDCr
+LtSTzIclW+FXclPRfQ/8Sh3cKLOwV8cxuXm5wUlSvKwkt2nwIhqkgm1sYU7zpB6/ZifFPUGL6x4
tjICh0QBryeHO5pOW5szj2AWNUPpjitpSHQfe51ph+LlXzwGvpZNpCkYcP7kfrSrAt0E4H4jPAej
AEAiF8JxsLc6zBFZ+1yTFhDBYXefC1OAZqUAfKocAH5VYvUu1Pift154m9M2M7Is1FQJS0vLrZXO
6Imku9duOQ21IPMSW4zHrF7VJqnIEw8rXwEK/qNgCJ0U46TxLcbltuTNAvPAxPxA39OExKyvbhUo
0yu6AHO755ABgps/AwUOd/dYZAI5GpdTc7IvHtX/A+kaTkPiBTxCH7Dm3EKlZg75+vdhAjb4Blz2
y2najsNc+NxCJwL54bgnDqqdGLTzN69zueICyBgOQBpAXUyrN7sUoCvlc95cFoeqG05PKW920X2/
EAkGpsVsEYfUVk2Z3ZZl2hOcHgaodMuPcVN1dwZrONkCcGAXvYKziXkvif6J5HR0bauXTicWFsNw
jVIwUyBjoBKFjVi7vayf8WiwA4PVvZp7cWvbNcOjLKbCQ02E5nNVX71u+Ey4yOgfpDPCia7vnqzY
tiZX7tSDHG5SEPCbK22ovO7aZSonzsnwVqaRlg2vubrh/4PzVgpLfnJJC4SIpFXPypquNMbeLgFw
rAyP4Ejbrgi3gjxXYgXN2srYNUUS7Er+uTuL9tzMJKAREnE8fFZI/Zv4t4FbgYcouLTnre0V0XjL
IQIbogKweTBWO3TxqbRucOuC+s+mMahVYrO88UM5rpD7kiOlvrqmsf4DlovTxp2AGbvm7bFRaw9w
kqyP86KN3dV/Q72Qq7u5emOWpeYihSEoe3MqyuCrvQNtd3cuRnh/zSYrQUHE/zo/3YLvKN/xYA0k
5QQb6nt85swlrJph8KtZeH9ykJfj1rOeu8os0PPZstekvFlbNIISRTBF0Z+9BM3A7URGaI6Hds0Q
4jF6iIOel8L1+WgXjKWomEU6d/KQAqdRWBwqdbEt1fr9KbiO1/SDH8WvJighBcym2VBDBImD8nej
lEl2fHdQZEMvYDSNeBtH/pD2H0eWNr096Ec/QkKNrNK1p7dphBs9CXhk1zyfJGzolyt+vLCqsoUX
lNfeq51onwTxxpm1NJRNCuy8MOM4uIJGc+Q6X81uAc3hm7by7vHalnmtUUfg5Kv9K0nbYDl6NMwe
VJ0v4+qhsG0yh/7jhmYBg1JaU8XHIkXmYmiYj0A4GS1eYu3IKtdppIUuKklOor0nCebLN0zNe5fR
3WE+9ANk/EzxBn/220h0E+gdzx3bwZvc03z3uCRSjjJe8nUpFpCrQ0D9V5S3XWAMgw5JL/aWD4a2
NCYsij521Y859s5Zz/pieUNdqt+I7QE8hVPqAf6CaweGseZFCaGfbcTVtlrgTNJRrNC+Cx/Fhljr
i1BpKvb5z0Tgj5YWr5sOKMrTU4QdrBKiat4r5ja3lRMSK4i2I23w0BIniG9lTY8D+xDZ48rvkdlZ
pI7eH87RCUZ/UTxrd9in50Or7lFeuN0N3CVQeIx6ShpKNSDhJyzJ16ZX+yhRGWUL7uSZmD5bnlVS
uIbqbzPuHptNwJyajxcTuHqappKOpkMwA+DY3z8n+XRXKz21VkCASw1vq+OOgDAIiObrPNIjsLhJ
oUAG8SAQgXT+eNd/+bncSO2HAklagG9wtICXd28pVxbScnE/1lapVZEdQHBD7a79abOC3AoAJuRq
eG44fgn6G43vLR8GnR4MaBQpumkd97IT7zc6nW1djlBxvsNFR3exrQfSTlm+E1pePcg0oQVW/j2K
c5uAYBIDvpd0h7JwqD1nB9pgy7V9FlJt4/V+Uq+stb8jadikai9c1iI0NbG8AdWKI132i1sQ+WD6
/1KcJfhZ0/OIJ8kJ8QcFppcNitjj+PpJaM6+6Zs11tgq0PzJLsW+TKK53Ck4e1EGOfHtdMcf3bsJ
m466oR17YqAGQ+ojAWOdBbx8MW/DGTPB5cmF7NoqkqmICR+usOCSVe8Uw2ZvoaZxPaW6L3kkMazM
CKh0V0wvHtcnki297ZBtxShrUd6F1/lY+VG9mhRr4JzRrP46oZGM58kNhvEYuWUJxsB/xE2qVHqk
SJTAoaSCRxxGtR3PJfQ3FCl/cDapi91UZWpE3D2IehT7EnOHyzBkipbrki1DgAczywcUNhPvuU8Z
n3497bm48901F3PSd4WllBN9Cc3yhenQw2GT/YjARijT6P22jFntUA50khiLFUuvr/C3Hr9d3YbB
pAfEvywm07rNAYUh8rdDYDyCtnIuSuvoUZRwJttqUHrvWfYsyxk5W41Mo7LJqCDHAyWV5H4dF7yc
n7uxrnRDwgMZDEgpsh2i0PIDgFfeDenjO/vGzWtQbtGxvayJlSyo4teSOsiJJ5qBq3uUT0++zSOE
NIXI+1EyrmVJwL5/eFERJ9F/izrFf1in3sJkMhw5/himxoA6l/03gdIK2goZTrawq+OGKoS+9h8e
oxmaX0chK7ZRxy57kvif2XUIbSAkEf+L1q23allkAxyjnIAO5UwgLXLUKhpQnBPAhQ/1A3rVHgii
wzrW7IFuQktvI96ol5hT0ffuwuJ07Cf624K+/lftTe3xsbkx30PRGF9ZlDz4kMTfDFzP/Hbjgd5t
lTUPA1JvfDQzzZCgicU/LGU+BehWlRuGiorWsyOLgYuAYEbtt8RfSgt2tjilC5OpFDaeWe5GJuen
P3UacOFl7XtIbSo28Od3vLTyikpJKukGIT3xBZuceH9s58wkHq1jMl2OUe7HvvDae1YuvwvSWmc+
VToDOAj+cQUCVw9PUbEHmp8NqBsoISONtIYw/ecJuanVeCgy4JIRxWqrsfU/VUjBMU2af74DU5fT
2ZIEkrcfX9rx/OlX6IglVKu7bpmj/pS3Cu/LVYmtLWCx5tasDLN2aauQiJ6VEPUzP5Ei/pb3AMa2
Fi3vMgKP1B6drl84J++rCQ2QIGBYekzswyaO2Du4eb5aiChdjD66cPJuFP2/uRWPcp74DYzIsF2t
CpiH+EWiodFV5mmwg+B8opaVmT9EC2YulsMzWKnAOJaept0jiDabjHXLfZbD2Z4m9sg5eoun8/R+
s0kvCwILwvpZ4XNYd0fej6zPxil8S9YdzjZ3hRjc00XC2Kjp+unkVMRSOcFPDX3tG+uI4+R2Dgs6
RjjPvP04153TLP6BrlF6Sx64BHqX59T+IsAG64vPIYxgCb9ma72HkNUDZP9BbpdrxsA3v5haM1fV
SanPb9/sZLpC02MR5vsEVic41VFH5YGTaT6icEUmuyf1r9PWHc37nGjRuMHa47pkl1J/Ky9J1m3v
HWKtPNV9GwWgsBTqMMPwhfD4AdqP1SNplhf2YVGN3MT8T/a7T4Gn44xsV6mQCd/ZispWN6U1VKO5
x0yJlc1XOcfE8xspessAPnsxPBAV5g3ktpjAvjc118wdqigMThQGETuxoFxw3oh5tzNu2fA/53b9
s+SMcNenOiaSns3ckn3ZYmJUSOAayVsynIy9xQJqazMmbBbfKIRwvIV90VoaueSYOyKvBT21S4Wb
2BNTSrgetMzuz0dwdUas9YIOk4roE1MxgcioShcRwX5kvaqY7FdtJB23vUFn3qqLqmEemVjj5vPM
Fig0A4jnnZAd8myTueTB3yyNHZpsrozqqiR/FG9yZFfjEm8uSgtU4iby68aOO5rYWZDud0lfZkDB
eltSNWq+p1H5egBsf6bYgKY08F/zSAQrWgcQ2vOEqA9zQ0wVQLJ85IcRdyaVErdd1ZrzzwC81TC7
xsnr6laSa7Gx/D1FPSfacuTMs2QANO4MpIVzd8LLY35xjSFp0sX4k5s/FeBMLlYpbYywPysV5uhQ
kHaJUeGtKIKbc1R0CcSOVETmpdXwTsKo4mK/iojSW8AFlp4gMmAUDQfHQoT6Wm77S78drjMPZMOS
BKXBU7xgdMaAyQM8YCLp9UWSvLzIF5mwiXiCiZTeENhxE54Qi4mjFXjBOeZuRJfmBn2J8krEYMA0
j2UBQGDInfcJC+XwNSTDTuL89OWNGzJyPZVtvwMAYD3lzY6zae0QPTPD0NAbQ6XRdb/8xNXZIdGu
tWdun61I/2r4ZgB80lDQLvZ2oCPWgOYcPHdtt1EutA8/4iKdpDQGtZiHFA3OI3K1jkyrUAr+a1nT
+Y21shcjTMAXGL31JpFWchascXHpTqd5f0ZksRy3PQM5sM2Af0Xqq4B2fRdQcAOrQC/hLK6rKPAb
fFml5X7rPox3SSGoatS23OV0idJQEfRkuq1247muN9wFHdeCUIDqWlSmDw9xgOHFbXGYjTyd4WaC
CdyJet8eYBfKLtYMQgfuIQLXi9sXBJf7VpmscAwrNWORNr6a4EXIkvvZJOOD6FBuBN9gkQt009tk
DXVk+8m9A2zr1ZWSZeZaPwZphiMG4n5uBTE1QNCMcKqmk7VGQWJqvmH4++hwWgWKqcUbx5keOrxd
l1DNMssQ03cNT/V8kFAY0Hh4vOXtN4f1m6Ql3yMikuUznEKYDj0636WoaRDOHmUGHB2sjBkorRod
EdzZfWwcTpBZp0Z4A3f7MixXeC9Oqo2vhKbMcJV78CzfIe6mc0sOc++iLcBlCGDcKe6Rg7e9vJD6
6Bax1PHbCvfFQ7FdH+U51CXxH1bPXYcTPEu/R/dIHPoBotpEb/cT2kfFISczCHV/3CClw2OE31j5
KDJ5m+y8h54EGnGcC9mOIvPNIBKqLjsGFlDyR4e1lPf7nyW1Y6ZRUBqXfSJ3Mk6w+DDZE19k0wTz
n3P229vCHKmAhW1a9o+/FntCK8DZkZ8PDEJLBggVitX0C3mp75IuFWncDbiuYVU3rsb1UEHKS3nR
iEDwfsRpO0ZoKBHKTXQ84exkVp8/Oo05wyEwgwU+DO6gzUB/B90Ewa7X4kFHzyIkV/nAgRr8aI/v
r8TCH4jXKMzohU6vZ4jb6mL0oET1OOkaXftCKsNZyE1qAardf7yqenl1SoNYyjD6pD6QPhHQQUly
3b7XxFDyFa8erSeyHF9n1d1Df0QDrQ5dX+yqQwg9JaWeK/n5zu6ewWLX+zDdFUcZsLZ82N2mYAB/
FyEZYSp5E/yVRYR/X4FhniYAYUIPlLAFDOx4a291/NH8xv2DEljZVDXUqVrhtHsExTRlUpk8LRq+
7JVcsgNmmGxd2WUSk5P/YKrbH5JyZ7jQzXxrPN6rfLkIT5HGihxTnZ6KkM2Fy6Ek2+ZZ6cfmQfgA
NkIJ8M0Vnalfu7vmur7YIeOrnePu7XnJQdDCnjAxfH5zANLouwpfQTiAm4CO2HFyJCTOqbNzgzdV
2BmY4UuQDziWHnNXTincAG50hWWXqRIYUcjnzQeKw0jMgWnUsKf9oOi/lR9ORMGC5GPvCAuMJAAa
jf6uh5j4C9PfTgbiC8ywU/9wcmgy5yEBtMa65blkwZxvnBWp5mWZTCubPiG3Xgfpebvu9clXajRD
vZlAZN3lKz79huwVds1psdCVG5u95I1DAHYd5bPOtNIK8dMbP/L2MKmBA5gtLga+aeXvVdo+huv9
/IDNAUFqHQmSjhcSnsN1kvPCJ1PUrvesYb1pOFKkQGs3zypjUQhYs7xR2uKnilfrfiFM1ZtfcF3y
l742bekmTT2NB4+58RISzLsMZJsQQ17VOqZc5zkIsE5dwb1D22naN6oOjvxl8CRQQfOYKIg/jV7D
zLQhXPqGVn78Q++zvuv8HzdIZZFgtMoRGxW3mHT2d+0LL5OmEt48CQw12WnIi8/KxrsN3Vnub/Bl
sqSSk6Vrs4fjTLsB+lHI5MQmBE5HOJxhJKC9UTtyRqYxaun/wrHV2EovmvgZKu4qQKY0bBuco5/d
USgC8RWe410YV35M7ev4hDVIDq4RdUNpM8CtuvEdwbQ5cy4JDDfmv1khMYt/7qg8xQHV4Gkli0sy
UjSVXVqxJlPFylL8xsRwx6rlr2JhB2pvuknAPz98mTgIjlTD0ppZ05oEWbKqPc312kYmjbZirjKf
ljH6BJUshOzOcDKqdRHKYlov0LhT9ZiZUmDoYCNnX/UA1SU+wxRBYKjyKKWtEqFtMD4tWjPxJ1Ko
S66fSEAUWjL4Qd3q1R4vZ3Zgs9072ytr7T9uB7A0INDpZhDkO4QsDR+b3UcLYivR49a6tPYuOeG5
AP1BccnoKwm3OC6PURtTmTpZ7u/IrUMPuoW0clvC3aNLdjY9G+tJxlRIJ9N+KUIeedczI2m5A5NU
JKh1bA7PqwYEQt3YZYZk6qSXP6G51w+mtWvthKxRbONKDs1epmm0UpthqCdYmkSND0LfukBV9OpY
5V/FAQ/JXbB9jHFfsXV+zAaav6dXFYmXYwivsOqcp5pFkhzad0N6mzx0rriarJPxICexP7FOxUha
7GdXLDBsBXpLuPeJywMbVHgV+O0c8Oe9om8M8eKCVAjhZz1/qkqDozZFu6efvqIwO85MhqKKcc28
iRvNcD2dJOe9Z7wtwScXoNOj5QCLcifD+ZwW2LjmXuHz97A1intf5ayz+xM1edAjlCYOTizqkRpv
qTZM+R2ya5CoEExBIFvP9xdiYxZdG7D7C//Sr9220qgzuAdn9tJZOfEw4YEAJssmPm1Oxa0mJgP/
vv2FD1xAlO0v2wX7MWYie602bHHZO+F9tIjAe0LDXmGu6vwBD6pPCDD4W/6mQur3m4zH+ZzQ7yUy
DEB3d2CubSSTkCSa6ow6zzgzzhzBk7vpNFExMZAXInevyblPd6IFxhwqvcmem2oZJyYDB3B/PAFz
p2yKbaiIgXlv0lZExneRit73QbTc51BXUoLVUZ6Dhxlt/f1aLqFk88GvpaWlCExIrhKEXvCZzXFC
ZEN2lCMQAgfDt8NMHw73im1IBektJoN5IUrcmjSbSmXqqAIIq5XFfrxt8UnwYIzDuRcO+YAZgm1/
BIWlWARNiK6JVNeaOaxWZ99zDqnb0bj6tjQ+LAha8jFLjlTwr5fQa4w7k8Rddd6jn+E6IagT6wnq
oU+yChxAylJojsqfrjj/EldSdK+8JXy2BImJTBk8fpjm70VGiYDgmmxvGKbl+rOsf3HpnKJ5bnxY
KFXFjMtodj6W+95eIxon22IDOkdbtmOvbp4iSV75HojQBtIUYZ2/zCp6VJdAUswQeHwIOlv9Irga
hdI+7H7Bn0FIhepihH50e45WRVMm4ry7xAEimk2QQDW68OLjTQ26OGFVWTpeh4KLlTrvofi0Brab
f2Lo7pfvvI9kVgQOCTqJECtWaOH6UOW57gYVJ8wjJEOmHaW5Ik659GPTPGOOecFsvTjSMd23CEGM
ddP4lRg00ah4aotxiSeSIrIwSFglmXqqLRX/vdsyZxVYgpYxRG71wzTmre1LX0psKYMz7AwX9aiS
nXrbAWVv3GcHXnlskD7AnUfCAyNYEu37IB3ewXM5wX94iK1D/xxZVbVCHsyzSwJOGQRnVuM7gx5J
LVJFwSoDMLj7ESpjHd4Zu0fQvMzvwwyDWKNMSNueipR1qYeOfi14ve9muJLWBNRSX2rt/l9uUX0a
Xzn7HNsPWdarjPZ0GHiUkbqZD/9GyKaK6fScrSJv/mZrLlF38nRRFm+q3YCYxlvvS4ctbOlvM8DH
pPNU/gMUZCyN1xsmXqUaXwCmuzEDCwnSHoqdS2BdA2PIaBsSAsf1mg0V8sVr/J9HC+FCw9rhJIvY
2xlQy4Fq7n78rrxG4yq0P1zdH03fDwUDqp7i8KTByBe1ioUiQ3gMIFu+YvVSwG4a1O9fgw4Hm0bb
f2b4y6JeEFFDaQewMmly3jqNvxqgG7X3gzDWSR/vK31ON0m297MYOLgqjoT9VHxDKeUn4gtptXso
NS6QoOi/nOcEzhjqOi+KLPdBzNULBaQ1mikeNg3xgq3swCY5XwtrGGoQH55Zw8kTZMpYt9t+Lh2b
xlxOKuBvoCOUz1fbE44SDa8SRTa6wTtK+o8MjzrjTEIAVldQimyq2oqjqBUlGXLkQRzFr44+ynJi
tJifA5YL+R+w4lqcNYzH910U3sO3qXi1vEWqSRmnMt7FU1NULC0Fh62dMXBrytl7sy90WbTJl3Io
UO74edNZcMYyB5yemKsXfRpxLAY2YAgXy24xy8mw3HZuBRl9fN8mYySDgU2qyp7DLSVxP2h7DwOD
CsWDuXvxaczpTqdB6hKW6yjJP3GgHeH0WVrNqYwCjEi+vxEUW6yQKww7ES0E47zMQvGMraxzFQ35
vfQ5k9z2pDLyKki8Z/fcTzjywzcRtwb+9zjro9LQ7PsQ6sd7gB3AJWdbcA19qVoRjymaH0Hr8nJ7
dst7w9Dbe+Mts81btgLVZWiSS9YxeHChdy0S9uFWoLGUXpXfP8cZk9bgvR3PdZ6Cn4TWipU0xXSn
kC8T9/5Y3Rsdal1wTbKbOqMTqmZa9eXmG3OWoqYtfGA40EWwWELSTRz4Q0Gfj3iHqGsp26W6UHzw
+ZypJCuvS5pVXCkrCsdeiuB/YmJBRJrR7YZkIydiZsNoWplR1h2ChN/M233Sf6DO0xzhZGBuQSfO
11TfexSjVNoladWNqSAbRoF6iWlcKBHkr4BgKeQ075SMXsbD8NKA9mBxaWSp+M/Wy+4DRA9ExIqM
YzuUfT0BfYFs8uGa9M9LCKCLhA6PfBvuO9XuiKnStJR+5KfOSBQQ1g0whMOGWNgam4d2haAN2LeG
aqB0/ppll5/46CLuwbsOmWXKN91eAQFq4LxcpPm2oyccH5un3YWpm7FI8Fd6Y7WeUjL+odZZ4pr1
lROqF3KvkNqdne5MH0RmgLdZgG50udYTiPhpsvaVSateWxs39ZqJ8HYv7R2AeJX2d7YHZzS1A0Jg
Ukc6nkJO6cWwHlfRQtCdQbkoIVui0dcXzL4wbmLKQBRqimJ6nYFke/R0WjzaEJmHVh2xCZqU5GqU
qARCjYEtEzeBMmTUrhPO3zW6WOcpR5uudDSOMiYknG609pSUaUvOXmVJg9Yt/NC7ecLIBY8fO4Vo
+OYTijDcHgN57F/lt1X64KZyn8fMHKZYtVzaJCuTqqcKQlI1Hegy/QVt6hZQqMNMssEc25pv2PYo
NZcUoLoRBrejvfWxs/gVDy+z8LjOI7Nl5Wuyr6qTBx7Z5ZD126WHTnmDgIsSUYs1S0d9arLKSAXW
/z/L084CIBmGAGfTAASoc0KaKjiBSbHFzYZcH4tmsjTEnWBn+YbOCDkKkOiIJlR+06Il0RIvQfSx
BRQLDq0AthZZ+DOFivMu+93zKedIZ6k7/g3Lwu2dsMIMglng9FI9pFUaMKTTmPATnOEvINQpqcnD
X8H1Me3kBFEgUjYQEY+/nsigWU7bxx0qPdfhQhcSrg8DDn28tMmT9wHUxocFOoUmtrecdfr1+I/z
0IrWmL2Q4T4uurEa4lGRoAj1yPCAx9zrW8j72BsOSEa8u1+thlZfRRfDDyDMj4O6hD1/a1OI+NKK
fYtXE8jOOccqb2ITgcVfbt1pjFuaGbBfEsi9ZAMzA0sieXlkoNJZ1GC7nkhRqm309d6j2BXa2HaH
lcDxTh6pzzmJ1xR+2bgaEdHkkib4eNG8jYcdd0M757M7ESmTRKR0zQRxxxH28fnL+TfpqfuspgDx
jUcMHAQavx2q1yoBXKVLZEEyNnMmwRlTGo5xp+AwkVCgIezOq+qolehXSaM/ZWYFfZWvixrodCJI
qNlTaiNFa8ak2pRvLtWO0jmIOq3FCxhFuCg0v7ZpoVxGiCGeduwMklquxdzWtFg1vDW2a7Yhyk+2
PaZzdotxkwINGM7GQNsdjgOzP2rO0Pmog1yoeog2TfCKKHuBq0zm/i216VvzaekTERkebFM3fa98
vS+CXvDWPOeISW4Ao3mP5mqVGaNV5kVMrahIxjzq6JHjzj7lkJ8D0HW/pUZwSpyv+SBJWUSn1P34
gEgAXZPjepJSQz9ehAGBPWhh6gn7Qw8C73dJRziZS5DWXvuSDGZnxlr290yA2bJVZuBgp7+VWhEm
9F4iCHTSlxHj6F4jtNf+Q6TTFvTzgrq12zix5gvP8tYeqnA+HNiY7GKvxEuwo/7Xao1QpBQWQnvV
7rjzVz/XUQ2iwsnH9xyYZDtuXNNeWAx0qWKHUo5deCqkJ66//wx7btGwVeYqs5P8SpFq1iK46URu
VmwrKJA6rzMO6NzBJt+pkbIEgE0DVnzlZNh/EPt55nTRf4cnvggSe9ggCVjoClf+yaZmo+zZLfi5
qsX9/sTTDulK/i1iUVrADyTUVwiS9/wcawdXLXW2eP9pavZ0ysxMqPpdEdUHSsr8OcXPzsYd7TFK
N1KMBAWxqlL+GyY6tXfZ5mjFJ4zq5J3tBySNOa4tBNXTERpdQ48C5dNM9PYOfwQeYER+EJSYWRAM
0oIocBb2D0s982x8zlrUy3/PNm1kObD+99/lI3XShj+DJ3lOJiPb5P4MnD+u+85v0LOvCbk4aM/N
NUTUmRRkoW7o7TYBX+ENnm2Aq8kO4YwPuU5Up1/bcdDDrEx0G7afOwR/AgO01siOR5j3XmUy+SIO
m+L72/8pUDD0vB351GFLAjIgdFiwEgMjRuDHtLs96IStDqg5cEXLJsCMosMRXUAJGaASBYpgDtSH
tHlqOF/XUoKrwzDLi6/GKSEEuHD/QhM9GhmZ+UE++7KSPIBOwZOId8tn4qikJPIU821vFtodDipX
XI+4HjlyDdQfb8ynkdzp/Lg6eD7cVP2tGzW6Ikb9yImZU0bYacrgLFE6jgaDWoyRKYsZ7940XySX
RkhAMBa7ykF+dlwYbiqhv3zBA7vZWh8GBBkQYIncMnShLgqmiMkRmQOzrxEXPBU4Ni8UWaUQRUfX
SoARVq2aF5NQMMrgV9QbVDOlWVZQ46kCUj1qf34ZEW8CUro19Vxz9/s2iRWmltONtJQkBMdqWBeG
r2cW5mycxiLARuc82I+3zg40Etu8CpXtespteS0Qf8NntCGHiSmqwP83BJgDQL62UWn4em7xNdDN
zuipSRt29rVoX8sf5jYHqfD9EyA/uAP4CrXY/VtUTz5JAN2WMo0wbMzGygo5QON9ttDLDiHAqhPf
95hxPcmmDMiu/pBVdhs35KPTjwe03tog4z0fislrQj4DuKIGkia6plMaQfwFLwG4NpTt9iE3v2BR
emZuWyTqqcUzFcG3iJtCTvDE9g10TyPsN9L3UGPElYeeaoYEI/ZTlos/4uyqfz/yIbRJU6hzFbFG
ovBYHrt1JrezWWbk2uLEsiJeBBkzl34X8LibkphgS0iw0H077ALHW6nzqEzv1XKk9ByDFfSSVh1O
aCsyK0yMdGPqx8WZpXzEMLVGD20NgWhk914geJUyueSEx4ovomfUstUs9cb0Ym7xIMCBoVS/s91O
dKZKVx6z6bm/VVG43tKduqYZd+gJQSFQVV+DhL8J6SEQag7Dw2wfkZ8kYVlZWyGMV+zs5eqXAQyx
C8Mda1/dW8zruQ+4TbCcRCaG5U+Y4DnhAv3yb8D/i4yOECyCQynQILxCUvz58oEqGFX3KS9In3BY
SJlHbj1cStsfgOtnilhFRsZVAcOQTiTzBlZ3w9jXPtqcd2sAlOz7Vz/Zw5jBC4NIzz6GE0EiCvFP
SdFewnns/8nxs+pGWIiHcflPTQwXBZxtUkYuU/ACcH08ek1kaAYHbXbOMfrpmdZF75RZQSrW+qvm
BwG6zoz1ESJuaaCMrWABSUXAHlyRoi6senipEHGcv7Z08dCKUqZAiVndcpZI1cPaqFok3CyDKuKw
z3VNrdfoGUauVCQ8TB4eVbMe027Q7RffNOiUXyLSs1qGOJcvo9TxT6SmJmCo5qVoRB39kyHDIAWu
kMBNKnU4IVCSyj7I4iCigO7tByTAgTy5Knb9qiCPbB6fv1ALpfO6xi+OyZh4K/gZytfRDcM+0bt9
WkyMJ++RkiKRBGNw8LCLRGvqUoH66jMsm8Me9E1cu7YXU+Ya4xA6rg25KbM1w0j0XaGZhjeGRQXU
tbAl96zgXzpqWSC7uxBMNvRXUQRrKr4hXrTV84a+pIv4m79kibss5fOD5d0R18zJ5pJrL2iWCqvp
Uz2+C8eICnohNVtlRtgrY6D/eQ2nniu39wMSYjRmTZLcwETO5qqryHRQB/TNugrO8kCOSgQ49bb7
dJiMti6ftcs6TYmd1UJ9tJszkyUykd5/8Y1QDmIYcZs5/bl9WDs2Gpt/ZPTKE/OkETykCJp2XIIU
uaEDpMaehud81NOzs5li0pQ0RTDlfDLWzBZdU7bMMMCpUs5rbU/1A53h3qCC65X+rqqAlI3bMmwb
m7kW0y8xJ0WPN61b4AKJaakbym9CEcS88HU1aklW6pZ9lkIQSGcC2oHOk8zeU9BoQnPZu2NHtOfA
ihVVMHubApdrUKnw8T7ORGxOHFwhbTQ7uhO1gdCpkqYKMRkrTXOf0CDwqIXZFJ4+qCv50Rc+ywl9
pHwTi0INqU+9KcK80qqqEJ3+P3mU9r4YQGFsQpuv7yoeJEmkQqO1Tll9k4r/XpD4tnTwMskKkq8E
G+QYCUNVGRDnA4PD+zqhhD3PAkCJkqBq8QPQR078OI93/7QIgT+IFVkruVHd2otjVaffYahMX5WG
VnR8k1nnIXT/AgDWC8Tv7nzRW0lDOyC84ZOOmCEoxGJWIA3JWzzW0FNIAGLdznmUgWOI7+SxTmlL
PYHDUPW12VQtZLPOJMfUzg0bNnvLWKAvOKMhIchKcUy2g27zSf2woVEXD38zKDi/3PXAgjM3rkQq
ELWT4OF9VZj4CxYek0bdT3I31LQzDiuacaHvbfNiMwwNwI0V0R7xiHmbkjve0lIZUGs0j+po80Sy
a/dys9HA8EeRokgGu2DXjvRQkRmzssa3LrYsBjneABwQW+dgMJTc7DN/gJJjYZHKO0alIQ8w9YR0
iuiDMKhEwBiP1+TotuoaEKOhz/2xbMUtUmDSWwmi0pl+NMTf6snlfQAILL8kSwDu4XblywR3SZHh
JR9aM0Ks7sbm5tz003xLcxUA2tj9+5rlkKdLnb6xaSH4N2S3Hcb3+w1CKu4USSt/yJhzkafvV5NC
8tAor33M2drkIo0b/sO2SookiV44HR1Q5XWeUGaPNqA4ThWYJeUB8ZRFfs3JHlT1ysdQyzMU0fQv
NobXy6hPhx3p6eUUOQGouoGOxyCjIzAFZua66dn1h3DaCTE0OiYc3Cd9pSb0pd8ehXZuyz964LKW
Fs9J4cyRd+wLiq1Pl0K5geOy3VmYXMrwMEeOT7glSmstkhOyEoJLP1Pl7plIvGTzdN6/r6KV2tvr
Ax5Hs8B+HBlPTAQNlQVW0BD382VmUkdJfEn8iog5BXHueZiK+AzP7CijbFambGL2qzc/Bv++pp0T
GhvkoyDMlS8BEW0KlnLglfQ/UV0H9r/9udmcnnzsv6KAoYaa1CA7C5XEfiDgE+ULnbjHdHC7eSWR
M+yvoalJK+873w76xREqQUehJabZPiYJCQm/F+eaoPKxrqFiNTpskVzE4zii/2SIswdnRpS9KIL7
DY90r1ydlloTM46Efh45UkyRd065ziJDITji0XElJwPmjHmcy0e2ZCrjvN6sQSHgCvqG5MRUvBOn
dLhK3YHBLZPdYSWHCoN5LgPMTM4B9eDmPV7SHZnNU5p7Sjd43rTF6RH/kRhAr877XuOxgTX0YDIX
mNuoDmbArpssh56956UQ6oihPnmOmsmzjMaP2yzw66hWE2gRyx7znrbVH0fjl9lk5PxZStE4da4r
qcHQ1acOP8Fz5p9lbZFBeEkTdtKt8V8NJnO9xS+HNwB0ofKfTeOVtvEVKP8GnHO/KG10nB81kC8Q
vht5GdYglFv5pPEAFmxJxDsgnE6MEslx+l2FwQjCXHLRQMy1IIH2mC1CowU4vOXCGzsIAPLFix9K
f2ly81Wur4gaUp1UqQRKE4B7jdHdmVOvToMUB6Ui3ywBoZep1DxtVMTDFnDHJb3fXs2VGtgfSfEr
7khPKPT0zPdKtw1KL9nQZURjhCGhCGtgZGlaVYYFKNnS1NT3waIQREVKuATgE1U5sG5CkI9vJDfX
382LQC0YDJ9c6xRUOsYy4T/VaiR5yTkhb96NhvgzKdey5lerBqG1Uc/RZBE/lnY3IrFsFydQ41fl
aQ+kPr/A/awXrRF9FNfFdVqrVHYeG12GpdnANkNvpTCVflf5o3myh29WZSY2RUIZeiEejygqJKvA
3XIbAH0XwoR9r4ppE7cUMdNXdis0e6W2wVYFSVyVCZisQkhZpMnkWQ4DJknXOLbQpZcLVBuk6FAI
32LZlizt3HvtedCme2sdwPwBAUI4pxhZQO8nJjGDHAwM/7wQ40UYKWA3ReTZtmch5ofa3BBLWDOL
1UrKhxpaIzyUfu4Zx8qdzyQ0Sy9d8odKaJkGwndCu6YLtQ3LdUKVIZGcviyiJp4Xzqnq7Upm+hp1
4lsX3aU4DNiMxGpDnOgQ3wGo/r69iHGCWvtRhfNNOofR00AY1ln4jya7b+fHe0oavCeknBD9bK2D
NpYZkfzD8wHDaHU7IdHuVMb2rRhpQ9L6AaIbgX5CbG0/G9BXSt6GDu/Gwz2Oi6wj+yUl+bPE+R1Q
dNCT9yw6+Qef2tSHOZUX0WRq2vtTS/yfcTf2+ipUIzmrkepf1a/u+rORFzEL3JyHDotJq7jniPYM
nwfKDzY53hDLEmE2hRvZYUOWhkiuKayQ0x98nnGocQdaeyGuMRD3XJE7TW4urIri5HGs2+HMzZw9
RAA7bec8e7XgU/Bmpg+ILcHlyEYTBWrmraOZ+RUIpZZwTto1IH1a8TgwnZfw9JBJpPfMtdXsI5gS
ITsDLN9m3oSzALA3uhFPEZ2tReLXSEzHSIM30swYZDQ6O+7vgLx+WN/MfM9ADxnG877WfsqSWyfw
5HgjqY/jbgNEBMjpFDe1IXKQtUcpN9qwnHuvESFK2AiQVShA51QLc2v0nooIp3+EzILeqy8L7nQ1
XhAKlCcImCNkCg/3M22+093aTqt3aIyKJfla0gh88M7697cKlpfXydpkPcuh3KVxrYxKL/o12Mrz
ji5w+5axLcfooqnKyij95i7X+zjpNv7e94HjdqcMr6U8AaTLNy0Zp7ouFmYmEDxyCR4emetxGKsA
QK7CU7E78uGBp06m6Izz48lwLvElIegEfn4qfdjBxYvT3zSqiV+qApcDYS/UqmzQ6nVxf6KuQnBj
IhTTkTIp4itcLQZAPGawZHactC5vtQJtMkiM/W26uRK0t+ceJatOPXeqDIEmqnm2JT2FbWwFqA3A
y82+98ilvxm3Wz1SgtqpZB2LzR2QWeDbqVS85xzXbIJLUwGSsLqkyDw/vInJcYVtqZH+f2SX9qsl
qyIfx95xpn9K2Le5GoEt/18hTBIyY1dMVLe3ncnm2kzrMuOTQcoLNpuegiYBLk6SW+sxQFrLMI3w
bIfyTUhDhWQPXCMx7iOwD37pwXzJAUsF9A2oMD6fHQFjvNVOcc41X+sJdi0WBgUV428ThPoJI3sn
+Bv4ufCjagww3By236GsGtclp6SADYze6VeOjtsWd3023S3EDodoBxet2Iz5rlcdwkQje+qsDnEi
6olYWv5dCo1koLjgSGIHWprFL/QjprgWBIU/fIW1YelHcoukLraa8jlIqLkCSiAhzcaPJuwJyCu5
eNqs0kbB0CzXlE9G1d/OzRAlKqqtIc2LFmvNWDsMWlvme4EckR7FyjoS1iV4Pwgvk8ITzxk/CPpV
TgqYjB7C21MNP9KyBJBek7JkImxKFIixKMiG3lE5pUh+3Y0MW5VsUGGxaSLpIKzFF4/fj8wbVTsX
kiUlinhWvhfECpa4Th3sm2C5YAzkGpWDvYtfFuY5aB1i1PPet4tTz7DM9XlZrjC+YXPA8rRv8xj1
9WNadvOtx3MDTZfNMPrO1YhL7Z40jzjwWPUkdCE+OY/3luyy/CJyUFOixDDu7aJzeUpKz5IKDE0H
OzqD1FAWtcnT5CcCVGytf5DEKtNgni/S/e1D7t2Jh9WPXi4QxUF069lXcYoCG/NHQWxZY/YuWAM9
f/8CHd4mxA+fPlILYUw0uII8mBRiiUZyxeKgPKqbpR90rc+tp59otGL6Iir7Q5Xo8RO7ZjkcK3yp
HmAtoaTPXLMUeBNesGNgYYvBB3qwFGfSt5CvynNqsdQiJipcarZB+A+ICl4378WMlKGySumghkEX
TjPYjqUjtjn1HZ00c2fulZLhZWbM92UvdLZuNyK1xFpD0aog5sjnm9UlH8ipFqzn4aGLiRsyyr0T
CDguI3EXL2V1atxWheAsTN7Zoak6+tb2hE/wjGl818xa3uIbty9dgt9ajv94QJxl52UUbbKnv3OD
TWWtcciqb286YEIgaM6tEQl3miQQxEspkq/zdX6sJn/rbepOSQLEzzsmU+Ly15epK6MGFwjH5XaJ
VNNC9bIzNbNQBEEbwQ5jvkBpGUOfGB+Ygz0rSU0ujnePb9bRTY4Fq51BR1AQWagJ/zf2+vank2jx
2ThaKWZsh6l8YUO8vS7SEPJj/XYB5Hg0JgjMnNxzMlY9LBRG1W41n5eCtHeiTz212lwSWKKjQWZl
N7dIENtOKjjLYxURG0XlfSdKOHig3qGWTIzvZyy7A74IIhXuznrRze9RnmXRL84NDDRmf/pbjKBJ
Ludm7ET4anosVcEcN6EGLfag8st+O6OZ2/iCnXbBLDSm+ns0JlmuLSwlSJhUfx1hb0e9D5hQP73m
jNmLRXrAQGfFaqzYETEkqRVaMwARw3/NbNOdMiYSv9lr0RrCImKo+66FTIixpa6GT+KAEopkUuHz
70T9IgsRl8DULm5WUboQx5Ug7cvJ4Kul5Y7/JKp4BmlSvvilV13UJ8jHFLTqZID6XXly+u+90nsl
sY1rff4QmH4eS/w9OgVFUsCh6G8BVWwINC4camPReQsaNUtBiw2PxaclTQhSN8jjArw6vERil8+P
6oVNajqjEA+KKMQiTQFUQztJpWW03QO7U5ZszfbwIMMTJFeexTg8e1/VF2kyKslMpArd/C0lRi8P
8AVwJOj7d0Ha3r6HO7LOQI4V010YecC0dFmhbx2q7fa8VXjrz32dY88ZahEIllDrf0lY3s36M8kE
aPzw9UKgqrXO9u1AlYGyInaCxYvS2amNxiRPHI4gn5csb0Tbe51VuGV9MpX1MqO7EdvljHN5+501
H2NcTleoF+HKkGgWJR/V4K6B1lbwWny03c2xPA37jENNDT3goPEGwmrc5c9+3dpWRldh6JgjvNz3
+6+giEzoAztmxenyfSI5OFrGs0bxCJ68hkLuJzt/5is9plsOcU8hMxFj5oOzz9VY8+pILxReKeCa
IgKVILcFkDEqaDyg0X/wczX8uH4g0lHFAe1uE6H1JeufLp2Yt3AVUc/L3z0A/JfUEhIta/sIqGCt
qGVUqRHMt4idiRzSACnVOL7651y/Z9xpy8u3AywC/FSoIqBf/5f0ebfHZjLpk0YIZml/4ujZFYn0
SF89otldujXEzue7zOUa3xaVSF8xMpjO5VITz5gHrkd8P4YYcCy/Nzj4KKUPUcPVNZ1ZCVtqSvrM
CaHvkDYqI+z6LGV+/AIei2NztoHXaUO7H2tM3CQfta5RNF7UG5tmN/GCkzDE/+JUUXtNfLB8L98e
u7K6IULjq5kTyNuMi6Xho+GLffII0UOsbkze1SE56TffTMKHLhWLcYI2a7CNnR1qYlwmvWxh40MD
jeZDECytdGpp/aPoAMGK4DpJoUlp5OPPdf54uU3GIxJTzbduve6ID7nQvSuLWuTjalfPPLoPVMyD
Rjj9kIMFc10Yrqdc9N69oAI7rokya0RqsSD9x0CIFEICQrh/30qeL209BD2yE+/8ottElOXAXu3t
hHwz3BhhSUnUyNU636zawAq4Z5bPviQGAfIcuPs2KY1Slz/rUZuP+uD9CLR49K7MprPCD3YrizHL
+gIVekdIVytUF39ZL1vZVNJX/sPBLBYz0V5qpP40Ul5ftJDeFIJ98tvoLPtCSJkVUFaj+DluITgS
hiL4U1OrI5JKbF7dcBiqyX3QzO1KRi1qQsACP2b48sJcm6gYjfQShUa4iv/25Yhw98lcwFA1LhGg
csQj6knJROTNRjUNbcG5p/vN1v0yuQoVayXPQAiUr/dIBuLClMcRhaG88M+xcl/z23jfLiIt23Q1
IOLstMHR0SnnjVbAnz2h9HSXIU2tEc9XjfrDb0yBZ0ElmFn5rOvwU9vqeOQh6XhZBjmb6YKonCKR
3jcV9NBCDfcu94cCJirju+LS3E5XdCg3djxyszZv7doHzg6FRv/dXD7yu2VDkzzhUfng7bdwddgt
o3+pBmo05uTa0+YfFNMK14N7NL+LkfQii69NTx23ch1SQNTZi1rQWp12H7sqOgiDvbCqEX66oSr+
hJRyWwtOF+lO54t+9FwM+p0cWjJ0hi+OUcURG2XDzoQlcLwOt7vjyiV9f1T25wSbimNo3cJqmIcG
P9BEKdJFeC63ds0n96GUnbQAgTkfiJd8LQVrbXPFqPw26SNjM4jPgKk2lvIM0lYOKx7UhBw/yBqo
BMKofTfBRnS9CHb3i3AvqYB1GaD5D9qtpk7LmryOiNRQ8u1HLqrVBpg8NB07quaIv/Rz64FnEXIC
I1OPEv4Icr2QH+2L+YfS5ikmaZTqpStqDK9m52RTvA/6zQ5ics6X1XGu0hyoV5WuToiVYH6gRvVy
lXjOrSaPPVFN9+Jv2zRMGxD119gvVxXXO/buJq7Xgpt5ehw+68DEC4KedRlmwXTjjUf5Dx0K2HX0
kQ7n67/O+ekvqrQmKeb+HPXkrummhoX/24oI+rwMGjRf64DhJLH3QuxhK5YcFODnMADgyq9se0PJ
rAf2Os2LQ4crexcHB690rBbuJUUJQwTvet/9z4YyMfFuI9+UKMpGj6esPfII/8nemz2kjtV9F1Si
GZOyAqXfNunDyr/dLqjoLUbwSxPBvGQnaXwAMEZQiZjJx2ed7mJ0wifQ6ZRtmskCZ/PPUoAukFux
/307+lVk/PV22PuQRHj4ffZbUzaUFelYYrAA19DbS5z93dbeE/v1KdAzm9B3ttn2P7Os9Et/aVmQ
gxvIGQtx0+InS2IcrIH3bOfLowuWVa0MuY8kXAi7ZGDQLAOTNDYM6n4MpVR/iF0jo4Hn+ii1muEo
i7XdRMwSvN4ilvxd19etE7wczYOB+AxkTGcO/rr+zobXgnMN8jMmm31Hrcm/cnKZO4/LRzJ3J5Gl
OA20CXPkqt8KiIdp5X78ydnBTP2erxj/SOezGg1F4knGs8Isme6swMv/SMx00rFWzV5fyugCX6PD
AGmm2PABfEgQ9G2i/iT8io8AFvKtZuKXYbNst9S0Hw1TAVY+9axEQSjRO7zRFKlxBOwYepUFQn72
2Hn3yZ6kXbZAHXGgIEsiic5AI2dPgIIeQZmrQ6RiKg4BDYdbxY9cKKwaGSn8da3gU1V5T2UsFjw9
AryLrKaoHrDNiW2TdYn/cMJnDP24J79Nx+EKiCbchQr/JOUpQ0+6GnEBrOYz5TK0PhPhZ9FPE9+M
1QFrVTfsq85CjXzEt/up4p/UAfk2/3bFCumC2Ca5eU90/R66iI7JUyzzQfcowPPNpxXXX/dTv+BZ
b7rJvuJStGkFo123t3jQHAPElQ2oQCuIN9/EkDoaREDDXZLI+qjBt5rg4FkoWHs0MEsnmqmyH5Tj
aUcmpGPKLL2PQZtQBG607ATJ8XzrSDZx1K4TzWLiz5rCJiZAeVyYpLzE8AidVVa7d77c+sTlt1hy
Ywpw7nd0B34u9SCwXO7mSfi9d8bdwgzkJjdOBv+G/Ml90uCwWGG8NJfev0gJkr3cmxBcoSAuM/YI
SCBoQhrAc/LNp8P9/DOU3ar97iNbxwNskzh3YTolgOK5KgyUEXqFXBU7i/U0U3I9D3sYmoPE724j
NdBxIsCVwB9CoK6NvBI7p5ascUAeH/j/Uc4HvR6ZqPP9tCuaVKiAVZDN0sry8iPVuITw5A/exA1r
OYAjxCFvZd7k6EPNGez76/3WFhlDua3D+8DDY0Vr4S7ixzMv01GuAG9A6fTqu+YxhZFuDKtdduTw
2zbBMC8Be9yYixXykcqppWiqjXWnq7oLIgq4OzBPr8xeLBMIf3J1jF0Nw7YIxhe4TJ0yYY9Xyg7X
gSoEfW4kCEWmHlablK/JvtE7fYxuSSBZ3jetquJI/L/SFP3IDHdxv29xEMaK2OhgqVTHlgSQOHAO
ZQ2xhaSaw+vCjfKMtKMSPMjlrKGCFjUjKIvM31UaHxm/cIm+QSg92V0eTJWdG7ZtE6C4YdSYT8xn
NFx4HBehlAv5TIQv3jxd5DUksnt2s4dJ8NTG4hl7g7ctf6aA/4ldJ1hcDatCp46+zBDxbVaWT4j6
etl4z+78e+3CCuCZh0piFxvMn9vcwV7btrmYhctV1rjtnPkmQChN1zDSwU4OsFXeFcgDEYjH4lYe
dhtMBDlKXrV97TWjpgj5s/qOiRr1mggyEZ5EqBmgj/a/JkXo6+ZRSbFwCjNJ+IGMAH78CsTxXKrq
Iul61dge4fNRJVxG7uiLXzQKkv0CRXZeuCJVS8kh1rFJnhtXhA9Kw4zJ6OBeVnRiRF//e65si7nZ
jJRmDu020Lg68DVGNz+ZCPd3qBsfX7fdQWoBDv6opyWaSAYxP604zTcUleUyZvC4e61Qm3g6GpU7
82dbXGMZ6pK6ARzGxKbPjVo6KoTLXzGV6Hvso5aq2nHrNsnV0mrWlL9MonvYk6IWEDg+EmtvPmHs
k6SxAKDFRPMaHTjjg9C8+kY9OqzwM2L1pgCj0zRUX5vciST4lQNy6qFmI0MQ/pV68EtbTbzWOibh
9u4+H25ZR/pel8TsmJMfFPhZ+hL1/ms0KYu0LU/GNBZZ5zQ6A1WJCGZFWyGsqSyPzFOeg2j7JbAV
EABtnmwMUQrC1TqzS4hu9s5cE3rzz5oIRN1JkPdAql/hJLc0673P/TpD/+sSDu8eNdQI9jRRUKrz
7Vvhm97OuGng+NZ5cDoJAK9aeRGh5zc9ywz56m+tySE5xGnGO8ITMZY9M8Bc5SUGbca7EWtF7ln/
gD6O3L25wo97wvrJJGtWJDAx0iw3clyhNH1e8chv3JV1lpbHdRT3KY2mhhIPMQdZj75eBh6LIKKP
VOUWCgmHKf9G4fVxGQdLUlfz54Vu94XVy6dTQs9aQ5VFz3N9yDBykUQa0KQdhNi8a1qRoFPQV54w
LbU9sNbyOu318fymvFrLYpEG/OcpwK1fcEpNwPhMh8IOIVKOxBuGiWDdoP/lGKBa0tfVDXNQkRje
5z9GL3PP23vACHqKqIbp6UgmS2OEbmuAtDJ0JSKgbR2oJbLIe5VIVWxlzuDYVm2ZSMEsb33dqjmB
0Jre6Y8Ob7aK1T/OEnq9YJIPpsIgbbN8fulX+RIunN9xupoB6Z2X359EI7YL4Q1yUkxqshKBP6/P
9Uph2xOBQiLbQABhao52rquzqNnsiWnCnaEfBBVKdREqWOyaWCMK87gAko0SGcLHT5X52TYYM+Jc
c0cKGtbmbtUYW81vMeFV2R8A59c4LWlxdqMW3DFBRbrdMtoqNL606y9yYYXt3UaJ7b/tyay94Aum
lvYN2ar0gMcWoO1wiI7aX7095Bhne6gojftxdRfORmJIMtmG7hQFvGtMVuB/xd1IAFkdt3M+ttRc
V4jkBdQNP7J5XUvsMVFgtRVLrMCQr5YRADeONVohMVNjEU7rJwqmht2KKgPYNHktH4m1uHq0ODOR
T3Zt4awg0yLz3yq0UrjY5GUb+WcF+Fth/F25nhZXNMHF6SCGf+woGLcO8D+9hjoULWUmboYSaIxw
wKze5ljnM1xqzUaydOb1cPkp6DDrsgp+t+RmNDO4v5euzBHDcJad8sD3gM4sx/bl8ZtDB8o50iVk
bQFBE2PLBb8NmT+eRLdMBVSHki8nqeiy3pOYZOEG1jA58VFzlA3eVXvH5aNsu2UoDt8xT0Nwt91U
KiMSdcOLal6xQc/9TJiBFNLEk6DtXOKhl7FIYW2QYO+ZaWJ2CS5zNRtElJ1h2P+IJ97Gikk08GtX
2P3gbFH/F0GHrRZByBZIzhzykEqgvldHiKzSHhhQpcOX1twmvBbipfg7wOAQd7JvOcCeGuzKC8iN
ibWRSFBvefrQTYJEP734/hAPHKW8eum1YD47YdCsQz00Otyw0QiqJbLBXKhvYMM3F+/nGPvKmvLq
ua269OoDqF6Zt6scm5tw46+5S8RbBSLK1UKvNJnrai9GPQe4H8a4o65uSGczqjSHBmXKb5IOAsMF
/avbwZDU4b0Bi0rofdiNkjFHRVmy+VcvAQdRxOjpfdywn2FhuY6TG7WeZ14Y7N7eFKBvH5k+mG0H
QSpdMGuaitTBpeCvQNS0NhPsodUwJzVAMdQjZRpvuUo8Ukx/K3Yc7rKGASJmbQyHZrjLTPEueGyl
YC0kPT6GeOqEjFPo5ABFLJU4mGPFBr7wfFVCkzihXwMARQBAcRC3qGru0k2qmXLpkscyaFg5dQ/7
7AKxcnAmUZKt8waUDqYTPF+M4uBwPdGav3hrj8lMtr+oQu0/ZuHFXVi83cVY1rrpzBj4sKU0a2wm
faDnhaWAFI8wUZ5Fmg+rui29VvTf8OP6+M/fH1FIvduubKowrxA1WMu0A0UpNT8IwWjpRbMI6G5v
djUPSnBH/czi4ZGD/Msd2ackKn5J+Nbr+rqdj4Nd3nPuS+/i1YBSlE//7/uNS4Fb5QtdcwJXW98L
bRSmfVENvH0F3uLLoKUGppTnpOHqxAhwydABaWqryVqSic0Vyxz1qBVXRt5QRdbS0FpGms17ggLd
erw0C0ZCuMPOAZSeGZWTM+I8Ok7NgYDr+PRUAtSPDbDft4+j2PIv9Bx91/YCGFcWHbNg7G5IDYit
45jdkKjhVaRayIX/Zj2Ah6LSW278UI7xbMpWFGta0P8YrlIPR0UN2GfAZIxNfkWq5mHgKTzKG7cS
Ywb9gkQnizAqcMKOubGrW0IRu84I69FwphzQYYhdkjbTlC3jabXdgh9dVFFoYYy2RFAX76Pq8Iyi
C29C7IWUNU9WxKkuL4uciuTZ+ylhyAqrGt8MMcTccaKpr2A+QEntMm3HCyQZzkwdP8HWTfCC6bKr
s1iRlTFZx9gO3GA8p5WrCRZJqau07rvfQPYY/dIQmz9k2ByBDi4PBHndRnIJaafCyWg6NTy3coFN
DaBENMWm8j5VYkGz+4XovisxzBeJhbJGsevRBb14SIYme/9pBL362gN2UOVvqwQEvLj1GYFGxlId
rfvDsfEz9PQUV7oxZHaj2uGQHMJXl5Zjf4qCjhsCV3IJogruRxG32S3BTpm/yY68iYNou0aQKcx3
L3sYnZAjVRNKCUTtqfZtXS4GvIjPBt0ge8dnjqGbkEHkzpgjDwua88gcChTZTkTzK4k2JKQNyEfO
DUvgHDMROU0dcScIBdA6Jqktyj/+bZlhXBaODuPa3Q5hl45CzCPCl0riiibS2eRyL4VHqFQ/kUIb
PldCZ4z4AYJW+NQi2lFpRDDOSM+Q2Qk+xGmOwgmsjhp5PN+b9zb82qJudxzd6d2mHK8m2J4a/gAT
w/9da9roirYACRkKT147E/dV4p40XjzwKmbJZNsl1qFyMX+cDyrLL7moK6DnP2jE9yZJk+qtWYk/
paKfoIU8eq3suqs/1jKFBzQiQ0RvF3SD3Z3px7wC2gTQyYon0RLg1V4d3qncxB2Z+wRHu3qrlsNd
CDTI69Ao+iR31eKP6Tr5hEyUy9HjZZBvHnyJ2YjjXvbeAWCKGzUwQnUGs9htwr96K4QSmDmHUbFO
aFCxZpSNw9QS6n4/dXKtJ7CeoJOAuv5v29mZzSiFsC92VDQVjneoprnUjOMB3D+9KnxhqoElROIA
SCcEt/Ow5gJa/TyscSqzC/Vf2zMbwrlPZoB2C0PvDdrluTT0AZo3iLQmzMXAMFGDF4jjqzNwvtfC
6aozSIe0uzu+GgzteVPWdRaVgutZzmRSVSsFljAvcplZJMx/uThpPblxhva0B1fSBc0Fp5GaQ5FR
qE+vmcgxS7dBZ4a+aJ1qjH3sFj67aRR7xqP7gECZMGNO93UkrfLDKom8us0Yc4v0w6z5UMUntWYQ
YbJK1H3xJqsQpmAFieW7SqeKrHlvLlh5xy/0hC3/GLze1J9PVA5Dw1dN05ChFczFj1jNyPGzAJtG
4IL9TckK11TMQwyubZfWLGh1Avw+zo8bNbna8TxxRNS+hIYn9GDp8E8m3rKUbX4+FiI7tuGcoRyk
yApgqXc7nbZuvF29Yz8xp/leHBeX4vdJXZ2yyOD2IfUBH+Vdr0V33TFo20H9K+uqz7LkbDRwDvbM
ImI8KrrYdifjRp+tZNOEpdN1Nn9BtXEs1EcP4eTcYTKMYYkarHqSHyBPascbSXcJj6DqlPz0ntVt
bY1alQR0Q+j7FH2MBd5fBouMqAUZf79NQ8mSNlUxX1gOpc7tjHsFWJcuDRjjYzu4OC8zUaSj29JT
4UB7PT7N8kJrhDRSMN8d2l6dAzNqcmJ5tYSGUbQ4h6RWxp3hNjovNtiSCHSyD71TT6M0xykrfL6t
YjbVPjiSMhWYGojGXPf1hQX23ORjpvpWL6d46nbXtQyFdH+xKIN9oN4+o1czn1XEzkgVtLrnyXkm
sPrddAz0qoBrY4HPOKzK7mMp5E2UVk0M0/dlMxRCVGCKpKiaaPRSQVSpwK9D9fH0/Ed5pcMOOYv0
QCUDzEpx4Dwsui1VG1UuA7Ib1EI3yczZmwA9kTWcHxO7hA9hyfws8f8ZYtxsiUJ9qvaSGX7X/Kx1
4kVS55+/GejgeN5DQ5LbBXqICcTqtcj/CF4nAziRe9P7pkydFUB62YXMT8ebOjLV7ni+mOdbuz9Q
/E9FlV+RYVK73MHjX27Vz9mcBvSRSu+8GZG6/PVfR4zdUC7wSzlc+LttmbhTtgKBatqgRW7HIvgf
Z3jn9VldS8uccTHYODkozC6URuf0sMJYgfpbxrbzGqiyouPIN5hbaQbOYX+AzWA7oPt4gjUMZ4ZE
hkhjfuzVG8OI1WYK+6TcMTL0jjuk2/FASqKgBhT+bfP0i2R3kHmH0Qc36jzrJvMUbD/PADkEFLmF
r3U4TqltNbR86pR3SUqcBfCzt8hHfP41dpyRWfZ+d5kCzb7SNtW2qu/f+eIcTRB45bwuYImrTO/m
bQFbHZ456pNNdJA4ySnahA/TckO5EUK/THrirxgKX1aMCWrfP7ZzmlY2ZNeTi/eprfA3qmwnNV2j
3zdA9nzt0ZMJqMfsUAcQA2HqXcCMHuawJYrkGtGO9zRfo6tLqO51vM0bEtOpTfvyxjBzojLDC+V0
xWxNmDHRgJ8Ng0nFQDGUVoVcCHcy54c0ApIiRoWaNZBb2TqFjYmjOe1LU143AgrOrJYBGQShyomm
dFTGppO64r5VEJwSe5MnL46NVLWoVx4qWiiIPPo8y1RPnut99SQo7V2baUbdcRJ4UftyVKt6ViWd
8uB8MaAbb8XtPBt2z5h4HtKk0RzTf5oucw2sFrlrAmNC22N2Yw5R+yHQkjovSZjEG8GetvfJQ2KF
LvL+aYgiPRCNekhcxS1TlXiJIYQhALUpGWq2IFfdsbraxCBpTwWRCnfwmwIRkJL4Sn3hobZMEzd3
l/e0v1Zyqxlyh1CHGeYX/qehgw8riRt4bRovcauNCk1I5MZ4UTPnAFPKrWmva7FqcUme7kK/C1DT
E510btODJNOzbkfxvhwvGXzFT1aQSZbJg3wzdmM2iwqYqIfu+FE99bd/mHeEuqQxkBAe4klVcdof
sXtSQdgPXkbfXUEtvoeg5kPhLzd5MzbnEQnlkOUProwwaEYNdrp2OCwdZ515Oz0C3iDN9qXHqOOA
1YXx0ZJrn4e9pM2VWjy+5IvNKOpt5yVkdYu6UilfTak+wTsYsZ1MVqqk5wACprBUAlGL/KxXrTDv
zj3OjwtMEhcrtH5EpBu9cTnNM9gQFFBLDspYNJCiuW8g14GBZrKkbgvpDYXUKjQDMacLQ87y3uCe
8pnEi3XM/txUKukEx1xQ6lz5XbPsFh+KalMvnE5hcgN3vObebIIYuO0GEvtVWfr9kM+w5EoRNCxn
ycrxNjVhVpJNLs0pHGMYa7EqAMMELxTxGyG5r4dq0wYcuGuy5P1Irl4Qow8Z9XaNwhcmeCSd4Zkz
NrAjoK+bGIWYpEyizCJKJU95dIF648A0maqBrZ6KX4B3tmDu01lwazbF7T4vNY6K54Oe5peOecQp
ULBCnmL+O+n5w50hhJ9AACFUWY0sLS+12fzGKoHpTTALHwo2dZx3vtHv4gK4Yf7g4h2qNDDh7xeJ
ZvAiySzHiwkoaR21T5XjNF8dJ6/qIYSysFX4Bqu5/IwPBmRnnyZvhgx2fbug/NvVbkO9Em0/VTMf
znmEsw8CA1ajiWBMvY8dRR15wupC06seNkBEu4vnQkTjfKj05jSj/XzhOhRMjYt0B3xcUs5upqeO
3TPYgZAg+Oh+zuFyDQp8sXiF3R/7iXuH8QTXg50H/1n8LDIWiikkECE9cWOqcIt/am3FlgyCiGKs
7oT85UcweZkNrM02z3BD2y9JFvw3jt8V01R33/ZBflY50+6tHXJOJeCuX/eUXjjmrXPaIO/Kxjkx
VMt6ZSsd++WSpcH4+Yfl5NLeA3Hs/H7FLuDigiih9hhh3bui9iLmVI2t4ZnqA/2qRYFIQXVgf93j
Puu1ZvqeFlAvi3BpS0sxqO1dCsGcoDn4VGrh0VMMtQD1NVuqAdgyBZ/vXHHkmmK3D5H+oDvRXA7Z
drZS7Q48BvjSdinJ39IlkTNV7F4Bd4GVFHj5Q5biEog0U5aLTG5/mdPQyjl/uPHlsZ28rOKoMt5S
jeiuC3OAy/NIALdKTYRQmqRflf3QsejmVNTdymUWl3TLnR29y7JDuU76XvdBRIWiDHOBzaOH3fSj
cuYBKzgnyniKXFbiDCLUJfN5Cns5Vbxyuay2GMN5q9FPsh5GWRpeeHt06gWbLNgCUX8SUCqUPljK
sxdZHN+oymgn/1W1izGFve3kmHMMrucMDWCiSfSjOcnr3hDcEug/9gDNWg8ho7DmQp4cJ0tpdOZG
GSCxXY8t9MNrJ2caECKEq65MjB91T8tg706BZ+386Ag6lEfhv0xI/oAbEex/woG6KjsshzwDziHv
Ald/lNnxxJHoOG5e4AH3K7mdaGwUfi6pv4OQMalsdeP2DqhmXu8KxIGUUrRS//FGZgyAjrFsSL1s
m7Gmuyzver19EW2t5vjv7jIuZnB2eYLvCgXm8tT52e+U2wKzcmtRdRJZSIc64KQsaFWJnlJOSuOk
O2UpS78/l5+FRs7bdH0Iac7/hrnRnrL7wCsKnH7NthgNo3cgassK/hks1YJUa/rshENt/oxSZ5mR
O7vlSyylwITIzPzy1CclmLb2CMObawQliBcPSlQn8kd7peFqND+/I4nTGMQrSGGPYmoko2WMuNbQ
sQAjVZ/TZHdpt65LEJbhuhUD0BGaW3+qtMhcmGsFxMidQrYLWnmh/upov5NPT0A8p4DACR7dyA6H
d6RYSFn0rJlIjXW3B05Bx+1bC2f4/kt97zuO7tgyk6a6o8xZErBdMa2RScAmUT3A3jgvwXxhD2uY
FgsiD3CICrpCkRMxJFXhqfsPFr5sggJLl5VRzA/hBt3j+g8l12S9x1hWILyN6aD3pb8x72tYHWmk
S6iuuWuZEp5o4k4hoVKYZMGIIevRwXEmzq3IjJZvHucbnHQ8RvUzled4VbqjIppQs1RuImUeYV7u
v6IqYxmS4EdHcEzAeKKDAWGEEs5FAxFtjS/KquOZ0qlrVKz+/HidnEWXC8a0xeag06i1YTbdZRBP
nvcz/ZfFxNdGUZVbKwAKe3tvtjVdm8V0Ib0iv4Dn/uLDzJfO6Duf5SP6UsfgomfojwmFyqm6MiM/
UcLVUDJIZ2Yed575KAJKltlHoWNOEU9P/sjeVsSxzNF9osjS7amFOo45VHavvU8gnO4stZl7X8vJ
njy8MAcdWUOa9oTMKW7F8NE81IT36bDT6kEGYbR4xyDTpWq5wSfalvdJm//13wOWOuPhGmzYGMsM
V5pfO43+we++CMZwnsd9P0cJGYJlEsNAFU6oKvNVJS7C9bpbxtbjxZgPJekoFMWjainGxj2wKvbm
NbAOoyodtGK7OS5ZZyzfHqZYkdyvMfr9fcd40T2c7KDy8tlzumfgYYAba7eXJETSd4H5HZO9Qe6s
Eb/R2YuGzpc/bzFlKwXfBLia9Nz8PBtkjuaJXWnV09dv9oWSPVq1B+fjdmrkIoXlHTAfexVtlASy
bhvcSn09XEzkK4mmvrqpUZK/S+kpK9gK133X+3EUqKTiq4IkW0W1UvzyeeP0vSmqc1Aq55pyceS0
gFKC9VZONnWQnk65XPMf8xGHpBStgrI59LS2um9x8Ld0NwlEUB1rwhDzolGGa8rBZrZ8D6TqZe/7
S0DE8oUAL6QS3vfa19S1tCko496DCM+rqUXkUptgo22+g322BFEfpCDTi6GP0uJXvLniEXUaIWeA
IkGKwamUOM+PoW7rALQnleuyOFXjyVbSqk8Qp9CJ3N4S8T3d7TgMndoqMq3r+4e0e0Y6KnZSaYef
efaNJRR27567nKLMt1MVSZxElVbll6p4jJ9DbBBmJxK4Uw8PAUn6r/ZJpM63ln8ItDIHLDfdbidX
cUrqq1KR7rpSJZxw3aD9teeLDFOTGTbCzOAEmmviE628/tTzuFh+Sty+dBrZ/IxtTwGOySwHhmof
y9JYUE5vlv8rOSKxy7rWa6DNDw/rzR0J9bTRFw5W87qZ4SpK8G1wQo2/BXpe0HNmK1tZ1ANXdq+z
FC94fdT1e57QfWUA1Pn8HUKGpIBkJDcjKKkKJidZSMWkrjPFDoqDhdlCDKqs0oTKA0j3N5aRrt0J
y8en3IyNlB51EmuIM1woNe+kkt2vLHkBOpTFdueQShIba7yzpNc1akzyO2gkeiXoPfM+Sj6GUESB
qbHcaGKUW0Bvc3B8+ubj+irjFqXLZLzEZpkziYt/HmfOHxewDlzpz5VP1GzUy0O3jZk0iNqqce9T
sVjzU/YSSgawf1DetqObJcDVFBvWp1/9+wfTSM81odn0pLicjVFkRjZsJtpR98ai2QGqtous8ttd
Q8bDE/0Qd8yICCMzRbARzx7kbL6j4tmmD87p+oX92SPa1ZzjfrsP1bUu7mPgQ2LwfUy5mDIlfaKk
T9MSgrmu38Nx2NFCflA2vl3+hh24EPxFvWWOEwHXHE1mUxBIv2gpxJlyRL2kRMqHVrVLa72LoWtb
SB/pWQ9quut7c9z7uFKLjdqwPapBZ0Eu4ugNnhzW8ywonYDYKkSw5RCeu1DK3L+NnE+nrTunx6Mh
x/d1ZEHJ7NqE+pmZQUYqBTusbiQYhKSdzhmFTUd/nZHsYI3RN5mx/kzR7qOJq0jYGd6QyDW2RIZH
J6H4RRAB7Buevoxy7DwSM6v4kmlLnxmWA4aXYCm5JBM08t7P7a+HOAV8XvOkrjnCHLlztoGbrS9I
MK0t0e0bXz82N0VhVxeWBiBWibbSdviOVLfQWDakqaV0TdjEzm9joWhrZG94me/T0nGhguibRl2k
ruRBWAxB/n/pxxDTjPHkTiLmXULvAipZinBLPaEg0k7iDnSpnS2P853X4oYif8O20NqdzvJax8QA
f9Uak0bLn9XxJXVjYM/YYZBMARc48scPlThQNnjP66yqswgp/9kx3ZsnT/NcaIR0zcaxoxTOi6dB
T/0XFb6qv2XkIY+B+lRfsZh5KGe6gcwWzzA8A8ioyxCnbXRhVjcECmFVeInw20N9US0ccCxayI9/
KhZO9dkdHHy79yc3+FwJMWmLTYiVG+KivUnCAEjtfxJ6y53e+FXlJTe72vqKdSPP1RjqGZitbDUQ
tJ6xhAAFHDQkJLlrA3vEMcWQvCYvZwEf2HX2ai++4E+VMRhR7LU/TXpsa6RIgR9UipWs73/sc9PC
jsPCVQa26cYGVUuylFnFwSoLFfwc08k1tTaSLUrUmEoaiLM80WpKL9feMsbuC09iwx8B/sJGgv3v
RuNLSsPM5Tm18QLHg5solgalC77AOONny+Il1yCiuhSsuAWuthcryx80dhAPBVrbWuhkanTb6MMU
rTQquJQ2/GzntEKYCGLmAiaHYKhlRp+JZQrYu4cO3di9TKmUD2NltmoJaLZkZqJjiyW9FDkO2luZ
Xu6inMGXLqO2bqfyWWewQlzRn+SIeheOel0gzj1EgSGoy3WqmeNjURzMxlhFz6dMKG8Pi/3ZzM32
mFNqgtLMVLt0Y9uzAFMkvovcAkPPPNQRm5WiLhPQzdX8AU7cmtrg05sJa8pnzFy6+MdNx5uYHntE
7QP/o3uPAX8r3PRXM93Z+i9qMjzX/JiJw3F96jaskBNF6mLgkYlhWesZahk1GmSeYOvj1Lfpz6Kg
V7JMY5pftqPPggWIPXOTnVQ/kDnwQeXXrBg9d9j1LIBoGKebmfFuPlbFr4S+zpqXhukFCwRiA8rk
2Fl+Rb6c4rXwfaMCfeHztOSVkTLGTZ+2pkUxvO9yOjfOOnvTEpakE4RlOuEn4Emqy8mwlw12zAdc
1QFv7Ds1vh82zNMzvNh5UxsOSp1Db0WzMCKf4y3XRQCuAoKnw4r5qFYl0nf3qa04fq1+a8s7Nwj5
15Kecc6JcRUihQZRcpXUjZzAa1qJmB0Tb+Gwy6PzqnChfs8e0GQMN6K3lZ3AbDhdHVlFLzcmGQsh
S6uaMSShYtOW9Be9G/HZ1OuW1VAwOLwNkXjwRmn2cbL3Dtk+u2hRxdlFpuCO1hL8IRmspzTod3qW
nlvtdfZKEDFB89Ih9rJwG3nqZWLY4JSrgybCkIfsriPkGXs0QSaeYXxlnygObgyuvnybFFHdep1w
rW6LOOOf8DkDedJBFkkw1fk4G0ZzoANHKZXzGPxg6DB3Kb1jaqbHO9i+29dP0hLhYprkESlt8ZwB
xw94gB6hHEQmY1E44vRacdjDMLwnTaaAMdwVRoR1SnPp7+cCweIQQ3zVzlv2JjpEjUs7wPCeDqAL
GWNUq5oSGmM0l/iDGAPn0Nyhk9o8tb1so7nGVF9x9gkiQeRdZkd8jo0r0R6nKHe9l/uScdmFMRTT
jl3AYJM6O+mk8o8OXFf11gjMGGXljrid93XsQ2u16IcEp3tHyrB6bq4FX3AY6azkxgd2smUADw37
dtDH65NXLbY1WnWRn5l177mpOadT/jcIbqNrUVJt+JsJzcGku/2Q/4bQeoo5f0osmeVuw+gIyPZq
wOoQVRgdh+znao5TWVzjoLwHgCfCXxfm5y/g38V3jHPN/t50aWGNyjGKKqCqowtk+FDHmK3mzqON
nQ6Y4Dj4QSTQmoF3UJHYV+9D10wHCgxRrjqdk0MohZouaZQd54Xx3eVpwuUfLTS+VXny479V2evY
bTN7N7jP/Kv9EECxkDMkJgUlWPmcqEfOy8hFH4Y5KF4VPiMt92uto1SERd4ryCOE9Yf9OoNWFSVw
Y8wLttcw45aRT4LGmteygbdfeI+Nfy/dhhguzvZ/bIFzByb4kuZ6CoP1omx6b/WAQsIo+XwR0hix
wsx4Yobs06QCA/gXC+ux81qc/b9usjqBQrpGI/+LsjWs8l7SlKDlt4AUa+xj2imhg2mLOrpUiOIK
t39raT3xqVwFDOt7TSgGHZavd4f6BJh45sQOe3NMLlGR/ycdy5pQdbyeHL5tlGB90oIj46wPFtLW
EQNCgVvNmCxiywd+Efuf+4A4qYjc0/RLTYRuOTxGnkmuvIWWwX4PzjVSEcz7qwrxgCaOgS8r+lFN
XVPFTdw3yy2R9sgUagzqeRiwFmganQAfndYznfmw6bI/ARcdtdx9WC99tXNNdLuus8VUyAAY/SOE
PwdPkchH+SplyGY0Kzywd9qqeGxpxA8aZRFYkHAbUbfeAThbHhomzW0emPDJ46FZGTi9qc4PBNHb
69NVbpmqx/mh5ZtQEPUqb991WGm8qHXL++FN3KRvbitUfL26WON34Gs4CLAfN8F8+Dk9Bx0JW15M
RpMiPUdn+3lM/iMU1NCfVDt382/M+P3qCAsv3/yMiTU3HOwVuIb4YNYAw6isQx8wL72+MEkcrilL
WYPDJQttRyn72bTz8OQDcywDslOoLtKQyPXIegawvl7UrXKdqz4K1ke8gDJ7G7vyEH8bz2t2kT2Q
Acsdv24Oez8mflTwGvEEa1R+Ml+/Z/8ynoyu+8AS7DCSgoxuFiG7Bs5geJDmy/nHd58paaaLavta
9CZx3mmfK2TzojLxAzxBaOpIPvsD2HOi1sodircGpBMtbNrgZTb/BnBomQfiwR5re4vHgv+fcvWq
sLf5EhO2NXnuHbp79nrECegpzwO4l0dClGRyo6iP004/Vu+kXEL7gQoQoX5D7MEyhXM0nVWUE0wB
TnG+Up4E3n76SKKiKWNh8UCZmAOwf3gF3I6zQgPM9/D25mF/S4N8Y2/F2tUnaoCLuCmSUQs0nKug
L2qlAv7ALQRNvTEj+Zla8UYhcH1dlSp9qeNcfWcbp9Mi6BXtBbl/Dz64tF2uuyb1TXzv4bHKrCkv
E8Rk3CKP/PnJxCHbb539CMd8wBki42M6dIkyBgZPgCgbu5lWaSEGzQQXFSXpIoy9XWukTLM05bpz
lLUKY4vz3FHorI87YOGnJSr/AkfDoLUrubrlU9flms0HSdwCmCx2GAUHcrOfIvHRqZxsXe2FdcdP
QX+Mdq+EcwdRv/f1ca4nn24dpEQxhjd0kzbw0jgM2GFTLUEWIpM2epBfvT2cJjIiDCpaBqExy9+c
kWS6aTAnyF6RClxVaEngm8eaFkhFZbbZ9oa+b84Ad5umwSUsJ2L0q7EX2SlrBlU/IORQePdoNZZ9
A+NR34kl0qcwWjFJ7P3EjIKhS4KyLUDjbjV8vHFq7q2XNK+sTIEMFb84B1PZbyf/A7ZpkDavlcoY
RlsSwVJkGvRW2A9zbFgGTAfmS6iv50JjJC17kD9DBgIjT9hTz4E55WBD7bUe9l9AXAsWS9cICyCT
Sno/btOrMxyW1w5t8yrphzLzoI14ct94DOoLluP56XsARo8CYnuocjPvnqfRgQZvxiLVXal1K6v9
ssdR8X8EdBg+bBIbJB2mj7so8Y4TPnNMv3h/T/TAXl/okGJHRZStVXJ1nhPrF4vXftHUmnuCAobK
vcyimk37/AeujXcsnm3YGEpDQ+xAqvefpmnVQ+kici+0z+fgTlhXpZML7twk6q+vEz9IkiT8YvQx
1FUX+k/PIo2rWnSuL5139aYNU80Ceee1kHQzir51ta8nKbs+Je0jQHjhILIoF1svp0lnIdYk2Siv
l5fQtNB/JIrgpsnGYRFw7TClgLJWytM020LpEnhrnUAZUHdN5V6IL0gEazIRN1tdADX5ND7ohWDF
HBahBm7OpCF4JJ89pz3LDS0vU7FMQmwVzL173Ad5kohNb8J7dH5nxLP64ZmDQcZoK6nqwkF5jf2k
zAZSziCF0RIoTaLPbblQfXtbbErV6gAaR37XgLpszeC/swOk/yw67z9chPEyAqEUZLJez6Er1/Mi
9QotVR66izUSu1axYbxH6rD3s1tm1Zc11UfyLaygTDSdqrDPzQ+hlLdb33Lh/zu7xXklibnkuzUd
f7nPFul96iRE0e/wSo+F4OrX/Evt/1NljHne+02vxgJrH4KmuA5Fh/WlaEIwa7kslCf1msmQxAoC
UC/LGVKfddWilG40xWldrE3ZhDgi6Y2PQIWraYrO307b19l1oDT0Y5MliJnAlbtWLc3l87qMz6Lv
Hy65z5Olw8sYd1ZD3DAYhDlWL1CsEyk+v62SC9h0PET8uDX3A16Ao8lP9W0Wms0mUDSFnLqTNPS7
b4z9gH952gOXPGVKu8FCW0dj1nlDartFSGUMLEzONrCDErNAD79mp+6HKtquRnLOXtycWcDEucYX
AUzZOst4CxoAbihXXbwSmCW8H9H9aHisYzYKRc6HRpl9STQKQ8tS/FX1N4B1dj0FYAOYcPxPn8B9
/xOHRiL1tJX9jtMh3YNUHcVyW8D0eMOBwfjXPkBF7f77lIM2KMurVnwvgsYC/JrTsnqQisRqmbCK
XqKAj+nE+7uluu76BGtEQdRGLAPDkj4salIVQyNrintcilIMEFTE5YPYgceYZ3FazmzAp11mg1Ny
B5uDePpVCK/Lcsw6wABoZsljll4Val9dHmqRyPK4ucn4GgxJEY5CUP9AStyGPoQgtC38ke+yQmVP
zncxP1DGIZorR4ToiIwt/PppSEFK1gIJJgQ7Ub01QLEc3WrbFHJdvnnaS3Vw+UfxwFe2lLXUO1Bp
U1V/87POPrBujqSXLtgAyglAIvzQIhY85i/SXm3hbJrCnmu298aMjYuvzUVL+XSD0wgasTg4aLt6
RNjTvn5UttzRbbjD2armNeW8G/fXBkzEqoD7/5PhdxyUNHc6vDjrCeDCQRJF6EjXZS68Q8RY8Q7l
AETdMinPkRwqP44A5hwpaLmyC7DI3b+98MsGCw9S4FJWU9ooBlu62kNxOnCwpaih8YOvCPZvq15Y
fZI3Ly9bbUXhl3qM9JACv3m58NVqvKTlt2i4krXB22stHA5+6QKOeBoV4l0MCwrDe/pTBjwSImJk
PoHZmvMjFOHTlNdx8K0PlERcPITX6Vcl9ppJA6dSNxOuCfEyIszVAT7iekHG0q0UpMnuHNQ96bb0
aBIQpwpJh+a/Me6KaZwSf26uKj7jP+CZIR7/LSi4GFCSYshVlpP18j/d5HwxnPeQRw/2/PFM+lKF
Lx3BnzauqV12vdyuRj0c5OQPLp566jC6V1+bYpJWMHjGLj4LrPoe100HUOu3HhWu70YSdVT03CFT
vi8N0iCSL0DVclLJ0b3Iz9Hinkk5h5bP+6ebaT4XlJswokVBdD8z94rpXSXdMH8bfq9XDlobcMq1
FLKxxWl42UpgHFtldyzkrtKZsjsSd1btzhFN59QIfzjIMUJ09ahOZ5J0q6RcIyjIO+RWFXRWtSxd
3iIQKNjVYf0/BRFzt5y369elh/SVT7b6fMpMLXc6M/hkVQlXIc4SNM/tFWSS1PZrlYZdJgtaG9dH
R/WLmHjImX0fpfYG0Gr8xCryRFI4H4syxZu6DLzCJi4XKpgcSMWiMiL9u2MmwQXqN3aCzWnPM72r
L4m2T0/TMp0xCRM7Oi3UpzFDGJI3sI8NQoi5i8t4xUvBl9rIERnSOFde1ohllW5P7Fi4wK6t9Nv4
kCl+kRF25Y60lQ9YL19tE6dhB/PKy6iTI/aOxDbonc2xoGhgbx14b1oaiN8B+WG4BZaI1FauU91X
YsCS3RO6bW4j9X+GTLuc3zf4xqc5N86aGYFBxX6CBP+sD1ikBLBrWE7J//eIf9JPlS/gbzuqLuAW
r6+BXpLDL2edxtIeFD9sV9+PQVxzz+YiMLH1Y8cTbr0Ur48VNRrvc/YMHse6MUxvLkSH5efy2CC5
h4paukVtMQneNLyeJVlJss5RV2u2+Wgo1iV5o1Uy+4kNAKMMWCAjwIrD9b6stsY0ijoh91Xd52FO
3VIo3cIN7+2eiBf1HeZX4kB0SIMBOGmMmgWuvGtmqu6/08rsugcl59m6XAE6uloKFqIVmd4g/dyU
kk3Buawee1JNWMdzhwc7XAofQp0PxyA3L+X7QWFK8qwxrVozCgTzTAp7RX8bDzMRgvcgf4v8AOnN
gUmU29G+PPABqZltE/GnMxqAEdepm50LkIlixhiXyQXUf/7Q/e1wCqUsR94Wt4jyETlh9fxD4VHi
dqeiTzT1CdAdxLNH2SGhcKYR0EuR4ZNI/OiE0iarpbUJAblTtlLH5gIpWXAOP3VyJ1im0PKX85xJ
AiMlcTgWHpa/02zTqLiZWYSiHRPGfff+Giv3oYgoguta2ShP3mfucLzh4zaUuWljTcLDSOoPATy9
EdaCxREZ32A3RUpI87ss5bqNMJ+rMm1aWsv9CnkhSGKfT4ArFISrrJezggK61Qv+P8uZZOZMz6rb
559EJ2/ap9vUMxCIX1Wj3T9rYGrN+FnDNL0AMea4T5Y8qB12eMMlcF32MfXM87sLWrMm+rKtH42M
M+m7gUMSnWDkXV3ZTTTL8gl3nCbrIadLxs70mtE7BqX6O1bfE1vJmp3fMxcYMWY8lm4+xAhVLkPP
jYBTlgwNX4lsaVBcj0gxGjLh1jxZdKWbmVkNLJcKhZs+hoxsWyJbftqELmUhf0mFxKESwO/fwWY9
R7bdambIgFY9/FKL5vUKF3qKGpkh2KseYpWoigUSgL9HIvNpqraIOZgD3B/9kp5yweuKnmVm1Ld/
UY2iaySOTseIoR2IKeDMILW+Fuhs4WLKpdn36Suhgqyh98yifmohAOchtasY9wimp63Y/8RTPzfc
ipSdvzQwWtNjYWkM0X6hA4UhM7Ur/4Z6haG89HaQVN/aUQeI1itScvqddyDDzG/zSJaaI04riHke
CdG7NrvIrINtJajY2lNGefVdjXyyadgr/FWq3GwbTEWTFJQKTX5H8iL6oFdsfsSeP9gsKqCmc9ll
bounIptUQmGJlXpP91DpQAXZwbPjKCgTDcsv/0yw0OQHLFP43KphPVQMmrKtZkX70FA/kMBvdu6F
VytmzEzrV1ZsTvJ5SNIdCHDHiU2Z+t6MvCYfqiNfazE79WJUPaRfemZThTOZsbbwxE9Whss30Bf8
5rbzgcQV2P4oIP2gATTZ7Qb5AiCDMpM/2/57DaYmDO6LO6NMEzv5ha29x1M89wvKoQmiuvS1KDax
Z+EW/oRovY3T6cgEAEGzmwwOhp/EhFnDFHzuFwW7KsJeHvYBHUaP54gbRaTMuKo6k1QV/OUS4gzy
fpcAXhGIjQCPmMz+/zEwk2hbktMhRcEgGNxml+3KHn+Oz46dhTcSvJ30rib6EvoK8EOh8eukqdFZ
Wv2DKYasZkwkCBvd4TngOW0WJSka2WG+YeV8xhRTzItMfDLOpkC0z0MEPmAQZuIgcfUtM2v4GDRp
B9IKqIRcutncoXYOJeT9oWOYkiOyiNhHoQb6LmFBHdqL8Xo1aVr8HYnn7KRca3gGFUOHzslZUZ1J
Jv3/+M0MTFcjbQX0tDtTStGmIs+09oxOjHkKaNn/LI0gpbTJLBlGVoFjdjHqyPHx+TKckvztvEgG
a2iWCmPvGnq5DzJ0Ay4d/n1GyM2++gwkzAhQUElJghL9b4MXhags+P6diACPZO3VFbmknqrYCMVZ
j2yQSKgNUsoNOVuGAhFJFhMYFIBG+Ha1x2p2X/L8/tg2SMv0LlPXgYSoOBCzhez8Zm6yOH2NcWxZ
gqJJNng8DGnm6J7R4sr4xhQ2NRegejQvRhIYssY9mbR1DTiW0bVL2lItNatt6GLx1rowlI66Z7FR
uR48AkBDGCPEwJa11zQzqIN3VGXXHaxkBotjc2qM33xGTonyeHBSBuSPUDHLNZfWrgZP9Su3tbQ/
IqN95TEofezU949cNETHhNxh6ZsfCKbKVALRuHzlC79rWLmCea0Hs9Q09AYgBaW5sYprcXwc2GPj
fZlDs7JNLflUwom7bxYBheqUyGNZ/tyzDbAPiOBD5rkh//7I+VQoa3lNlWcSbqV01yh3fH2tsfNT
Yd0OGAgtuQRfAChzRWB+azAM1kJTT11co57Sd3PwWYAG9+6Kt5TxMPvElEderIxHCESvgcP46VOb
FbGRp8oZmOANEZN5dD3LNeHPxV3E19orbvp2V6P3+tHAE0WlJjE5kDF0A8s463hkfftpaDS+4yQs
g38Xg+Jw93k8Ya3VrUYmm0yizFqLR21nUN/Zi+Zf9y4I5BjLqFaknaXhnX2zI2sfkYOcHw7D8HJI
z2Ckh3BkpRrqPUCt2DArO2MA2Ewlraz+Rq6pScvgqgl6pjjJTrCCHUaslMnMSzxPkHi2vcrK+pb6
MgqOS4rvo3/NFX3YtVVfsRK6Jp5SZCS9zhOlgm4RAn+Pteygqa+1X1wuj7mlUtN749iARMjyAT14
v+3jKj5XyTRg7/xtRI/BSTc4shkerLO9yKG+c9AQlNqJuWa/bCr7VXjP0HPgJYBAZb2fz0zpl9OP
KCiaWcT0RjhyOixhZAK8Pgvh+bPb6vajXWd5GHPlZLDk3XOzEgFUxzqHNmJOjNN3WWSPApNQS11P
qEN5QI9gecumYFm7MOZ9NjuKVXinlf8Yc7MFiUMlg3zolOuKywf0dxibOej/0/m3x4inL67eHNUk
nUZiezXZ1oRx2TcsdsA7QAX9BwQfw/+BHV51ctL7HiE5HtuIMMf19XZI6KERKThv6l0MsqSPFII8
axLNUAYj0NyVxluwBKWRxiGjTidmA1Br5PTiIHHR3u7hSD32eIifC1qfBs28No0Z6tTz+/ht0VPF
i80PnLwfrFnkRYBnWY+pkgUyPS6kW8XtMBKqkNA/anlThmQfYfyIOlDisrBOMHeCtS8LO3obpyKL
QulF9xdLflVhTdDMtkKO7zfjjKiha6nk3qtlDxB26WpuaKxrH11/7mLn3FK5sN//qyAFNWzspTD8
+UHVw3yqLMLMyHhwWoulRNcNf2Nk3tF2MN334NW0fl+C9tOmYp/nfeG/9qfK8FpmHXg2oGvP780h
reD9Ug6mwcb20e4lG5iZOZO6+/kLH+xRoIQsN9K/bV0MVlgCWe1oiHKxkcQuLZ/y8Ke976IYDurm
mjNg8RWzsjx7dUywIILJPm2uiTxLzt5DgqPwwRecMuxHsMVqhBEYFzNYEQ2pTgmBurVu5uYCSaVA
elQjZnVr7b0LhnJ2UFPwPFoImc06dZpYMkk2xEQLXKmoxILNXnqCWecHepbbv1OmM8xbUKWhdhmq
khoCsyIAuDHSAPnCRZG3zqr5hzp8rLJJoaXGUTYytJ4o2VNXvZ8HcDwPcVRsGFM84Zs8lW0bD9tQ
eI40Eq6xKLNcAnJi8G6YFjmrksrJEvC4/dtiDDv8s3+J4spDMY10FBdqAi4Uh5/NMCroGUCRlyqA
IOOqhg3IK8MQVtbxyclVIfLYwbkJX5ks57T4D0EMA+2T9r6hA+VYkPOip7zO2+e+kgzeZQf1uoZL
edCMGpJEBx4oE1xkTF1RUue4Q3vY+ORz0DCGjmTN5jLx1tYuHSkzPgc/W+CxQAVBsAXdeno063oZ
0YT+J7RZGYV/OAkuOU42sv80JA0A8nMhZvrwYVR5PiMKfugA4xnJZ8q8RmznZT38EfRdFVEJox9v
WKtFEF0FkX/37T8LWa+ikHf199A4nfDTJUSgOTOHcu9x0KlMww8dGZ3XlsifZVB4xW+KKYb1LJEx
80TawGn+vm71XN1+F58YCLy2r5vFKgLwj2mWu3ciAEkjzQfAARPexD1b66TsPkk3kJvwjTcy/z7j
lSNqaJ42LPXnOhJqNnaKCM+9HgrdxPBhzjBZfFY1ltCpvT1MKJEFGscyB+74k2mCknx8zFD0xEvv
JSktqMzmYkKthc0lwEZlzK76TpMJjeMlMQ2YS6pVVcQe0DaGRmJh5Joy/zYHITKCGJV/hHzhH6eA
CjkPLr+LKpspxBuy3PbJi61LMD44bcTqqVGGZcohl9n3dNSAhsMpiZrgFVR+cW2KqhBu68Ccf4wC
EsYdHVrr8XijJHo56Ere/p8VzpfD1V/MyHTbK8WA0K4CBVM0pS7jrktquK4LVPkjgI23jPKYrsKV
aubl1WfbkL1ObyX075TN3OaV3PQU5jxxcADDsJOoRt34/Wb8XxSZNT+HA+J0yQqpmZtpWWAbag6c
Mbmp1aVvBAuR2hC8hQFUrFM8u2A4tWkTHmUdw5SuMYWWwNK34bfoC0odEOEhT2qGWy9BhNtXOVfQ
G4w2Hm5XlktHpc0Cvj6cp5cfA1+6QHOPx1beSXGh+MZ2y/ysS0jE6qUzE024BGVuDgHcWX3/7BAo
17gnRTyvhg3P1/xzfjWYDeB6Ehq0LBR6fExdHW3LGCvv5HHe49ydoDrpcbz0RSqM7jps4HxNTNAL
zJMdgQuAchaWlqvHVOpD3/QMBqz9LwrEU72dz0Qw51UHCxlbUSDBqB54owltzEhJD5dcSDc+6kP4
p8Gpw2xL1TdwRD+Offr0x2k4nxDd0tsFJDdMkKhJlHxcO2oWftnz+HkwbNv6E28jxXRFyUo/mUdQ
cSAo2QDIe4d6Xa+CwxaH2Nd0T5bdfeyjzD5RpIlceTsUTh3HmwyP6tYTQWzDavb5k8pOIdO9YmX0
t0iaKOhuPpp9z0EaZu41XiqIaZVz90IUmVo8OA4QmnYjHvm/DxK4LuCwf4+WBlEYD7Rd9n/mOLI0
O/EnhsoQC39mNxzDcawBq+o8U87imEqCZe7sIQ+C9yWOcCdtM4wzQE5uAVEM9Uli+o3YNMauUWyg
hyvAQVey1qrFPXs0O7eWHP0Z9+DfAF/qts7LO+As+yTdXkyhXjFms9CwXo21OE0WZ4EaktPmvXaX
1gxLk24dBUo4CuuqEA+g8PkA4mMjDHAXqY5Jdq78Gb/3IVmbE45/9oJl7h9HAiCEi2Holg4IQpkG
MD8Y//LTwO/26ab8LWgBMB8OKNH3eq1ydc3fJ+Y6ErcsS45RhP5OKbGqrGIYjXC5IPtzfMCru6oQ
caxboK0V++8atDThTw6HPo3O2DK5ZVts77uusukth53CxAyjfXASZ46br8OxO1GchSdDk66PNOs/
h29IZZrudZ58kE79s1AFBUPirdFa4ZNl+XNbuy5mqN56HwZUVkys38CH9spUVFw=
`protect end_protected
